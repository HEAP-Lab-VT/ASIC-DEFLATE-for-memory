// Wrapper for the toplevel module, which is the combination of the chisel
// implementation for the codeword generator and the compressorOutput

module huffmanCompressorDecompressorWrapper(
         input clock,
         input reset,
         input start,
         input [7:0] dataIn [0:4095],
         output [14:0] currentBit,
         output [7:0] dataOut [0:4095],
         output [12:0] outputBytes,
	 input [12:0] compressionLimit,
         output finished
       );

huffmanCompressorDecompressor wrapped(
.clock(clock),
.reset(reset),
.io_compressionLimit(compressionLimit),
.io_start(start),
.io_currentBit_0(currentBit),
.io_outputBytes(outputBytes),
.io_finished(finished),
.io_dataIn_0(dataIn[0]),
.io_dataIn_1(dataIn[1]),
.io_dataIn_2(dataIn[2]),
.io_dataIn_3(dataIn[3]),
.io_dataIn_4(dataIn[4]),
.io_dataIn_5(dataIn[5]),
.io_dataIn_6(dataIn[6]),
.io_dataIn_7(dataIn[7]),
.io_dataIn_8(dataIn[8]),
.io_dataIn_9(dataIn[9]),
.io_dataIn_10(dataIn[10]),
.io_dataIn_11(dataIn[11]),
.io_dataIn_12(dataIn[12]),
.io_dataIn_13(dataIn[13]),
.io_dataIn_14(dataIn[14]),
.io_dataIn_15(dataIn[15]),
.io_dataIn_16(dataIn[16]),
.io_dataIn_17(dataIn[17]),
.io_dataIn_18(dataIn[18]),
.io_dataIn_19(dataIn[19]),
.io_dataIn_20(dataIn[20]),
.io_dataIn_21(dataIn[21]),
.io_dataIn_22(dataIn[22]),
.io_dataIn_23(dataIn[23]),
.io_dataIn_24(dataIn[24]),
.io_dataIn_25(dataIn[25]),
.io_dataIn_26(dataIn[26]),
.io_dataIn_27(dataIn[27]),
.io_dataIn_28(dataIn[28]),
.io_dataIn_29(dataIn[29]),
.io_dataIn_30(dataIn[30]),
.io_dataIn_31(dataIn[31]),
.io_dataIn_32(dataIn[32]),
.io_dataIn_33(dataIn[33]),
.io_dataIn_34(dataIn[34]),
.io_dataIn_35(dataIn[35]),
.io_dataIn_36(dataIn[36]),
.io_dataIn_37(dataIn[37]),
.io_dataIn_38(dataIn[38]),
.io_dataIn_39(dataIn[39]),
.io_dataIn_40(dataIn[40]),
.io_dataIn_41(dataIn[41]),
.io_dataIn_42(dataIn[42]),
.io_dataIn_43(dataIn[43]),
.io_dataIn_44(dataIn[44]),
.io_dataIn_45(dataIn[45]),
.io_dataIn_46(dataIn[46]),
.io_dataIn_47(dataIn[47]),
.io_dataIn_48(dataIn[48]),
.io_dataIn_49(dataIn[49]),
.io_dataIn_50(dataIn[50]),
.io_dataIn_51(dataIn[51]),
.io_dataIn_52(dataIn[52]),
.io_dataIn_53(dataIn[53]),
.io_dataIn_54(dataIn[54]),
.io_dataIn_55(dataIn[55]),
.io_dataIn_56(dataIn[56]),
.io_dataIn_57(dataIn[57]),
.io_dataIn_58(dataIn[58]),
.io_dataIn_59(dataIn[59]),
.io_dataIn_60(dataIn[60]),
.io_dataIn_61(dataIn[61]),
.io_dataIn_62(dataIn[62]),
.io_dataIn_63(dataIn[63]),
.io_dataIn_64(dataIn[64]),
.io_dataIn_65(dataIn[65]),
.io_dataIn_66(dataIn[66]),
.io_dataIn_67(dataIn[67]),
.io_dataIn_68(dataIn[68]),
.io_dataIn_69(dataIn[69]),
.io_dataIn_70(dataIn[70]),
.io_dataIn_71(dataIn[71]),
.io_dataIn_72(dataIn[72]),
.io_dataIn_73(dataIn[73]),
.io_dataIn_74(dataIn[74]),
.io_dataIn_75(dataIn[75]),
.io_dataIn_76(dataIn[76]),
.io_dataIn_77(dataIn[77]),
.io_dataIn_78(dataIn[78]),
.io_dataIn_79(dataIn[79]),
.io_dataIn_80(dataIn[80]),
.io_dataIn_81(dataIn[81]),
.io_dataIn_82(dataIn[82]),
.io_dataIn_83(dataIn[83]),
.io_dataIn_84(dataIn[84]),
.io_dataIn_85(dataIn[85]),
.io_dataIn_86(dataIn[86]),
.io_dataIn_87(dataIn[87]),
.io_dataIn_88(dataIn[88]),
.io_dataIn_89(dataIn[89]),
.io_dataIn_90(dataIn[90]),
.io_dataIn_91(dataIn[91]),
.io_dataIn_92(dataIn[92]),
.io_dataIn_93(dataIn[93]),
.io_dataIn_94(dataIn[94]),
.io_dataIn_95(dataIn[95]),
.io_dataIn_96(dataIn[96]),
.io_dataIn_97(dataIn[97]),
.io_dataIn_98(dataIn[98]),
.io_dataIn_99(dataIn[99]),
.io_dataIn_100(dataIn[100]),
.io_dataIn_101(dataIn[101]),
.io_dataIn_102(dataIn[102]),
.io_dataIn_103(dataIn[103]),
.io_dataIn_104(dataIn[104]),
.io_dataIn_105(dataIn[105]),
.io_dataIn_106(dataIn[106]),
.io_dataIn_107(dataIn[107]),
.io_dataIn_108(dataIn[108]),
.io_dataIn_109(dataIn[109]),
.io_dataIn_110(dataIn[110]),
.io_dataIn_111(dataIn[111]),
.io_dataIn_112(dataIn[112]),
.io_dataIn_113(dataIn[113]),
.io_dataIn_114(dataIn[114]),
.io_dataIn_115(dataIn[115]),
.io_dataIn_116(dataIn[116]),
.io_dataIn_117(dataIn[117]),
.io_dataIn_118(dataIn[118]),
.io_dataIn_119(dataIn[119]),
.io_dataIn_120(dataIn[120]),
.io_dataIn_121(dataIn[121]),
.io_dataIn_122(dataIn[122]),
.io_dataIn_123(dataIn[123]),
.io_dataIn_124(dataIn[124]),
.io_dataIn_125(dataIn[125]),
.io_dataIn_126(dataIn[126]),
.io_dataIn_127(dataIn[127]),
.io_dataIn_128(dataIn[128]),
.io_dataIn_129(dataIn[129]),
.io_dataIn_130(dataIn[130]),
.io_dataIn_131(dataIn[131]),
.io_dataIn_132(dataIn[132]),
.io_dataIn_133(dataIn[133]),
.io_dataIn_134(dataIn[134]),
.io_dataIn_135(dataIn[135]),
.io_dataIn_136(dataIn[136]),
.io_dataIn_137(dataIn[137]),
.io_dataIn_138(dataIn[138]),
.io_dataIn_139(dataIn[139]),
.io_dataIn_140(dataIn[140]),
.io_dataIn_141(dataIn[141]),
.io_dataIn_142(dataIn[142]),
.io_dataIn_143(dataIn[143]),
.io_dataIn_144(dataIn[144]),
.io_dataIn_145(dataIn[145]),
.io_dataIn_146(dataIn[146]),
.io_dataIn_147(dataIn[147]),
.io_dataIn_148(dataIn[148]),
.io_dataIn_149(dataIn[149]),
.io_dataIn_150(dataIn[150]),
.io_dataIn_151(dataIn[151]),
.io_dataIn_152(dataIn[152]),
.io_dataIn_153(dataIn[153]),
.io_dataIn_154(dataIn[154]),
.io_dataIn_155(dataIn[155]),
.io_dataIn_156(dataIn[156]),
.io_dataIn_157(dataIn[157]),
.io_dataIn_158(dataIn[158]),
.io_dataIn_159(dataIn[159]),
.io_dataIn_160(dataIn[160]),
.io_dataIn_161(dataIn[161]),
.io_dataIn_162(dataIn[162]),
.io_dataIn_163(dataIn[163]),
.io_dataIn_164(dataIn[164]),
.io_dataIn_165(dataIn[165]),
.io_dataIn_166(dataIn[166]),
.io_dataIn_167(dataIn[167]),
.io_dataIn_168(dataIn[168]),
.io_dataIn_169(dataIn[169]),
.io_dataIn_170(dataIn[170]),
.io_dataIn_171(dataIn[171]),
.io_dataIn_172(dataIn[172]),
.io_dataIn_173(dataIn[173]),
.io_dataIn_174(dataIn[174]),
.io_dataIn_175(dataIn[175]),
.io_dataIn_176(dataIn[176]),
.io_dataIn_177(dataIn[177]),
.io_dataIn_178(dataIn[178]),
.io_dataIn_179(dataIn[179]),
.io_dataIn_180(dataIn[180]),
.io_dataIn_181(dataIn[181]),
.io_dataIn_182(dataIn[182]),
.io_dataIn_183(dataIn[183]),
.io_dataIn_184(dataIn[184]),
.io_dataIn_185(dataIn[185]),
.io_dataIn_186(dataIn[186]),
.io_dataIn_187(dataIn[187]),
.io_dataIn_188(dataIn[188]),
.io_dataIn_189(dataIn[189]),
.io_dataIn_190(dataIn[190]),
.io_dataIn_191(dataIn[191]),
.io_dataIn_192(dataIn[192]),
.io_dataIn_193(dataIn[193]),
.io_dataIn_194(dataIn[194]),
.io_dataIn_195(dataIn[195]),
.io_dataIn_196(dataIn[196]),
.io_dataIn_197(dataIn[197]),
.io_dataIn_198(dataIn[198]),
.io_dataIn_199(dataIn[199]),
.io_dataIn_200(dataIn[200]),
.io_dataIn_201(dataIn[201]),
.io_dataIn_202(dataIn[202]),
.io_dataIn_203(dataIn[203]),
.io_dataIn_204(dataIn[204]),
.io_dataIn_205(dataIn[205]),
.io_dataIn_206(dataIn[206]),
.io_dataIn_207(dataIn[207]),
.io_dataIn_208(dataIn[208]),
.io_dataIn_209(dataIn[209]),
.io_dataIn_210(dataIn[210]),
.io_dataIn_211(dataIn[211]),
.io_dataIn_212(dataIn[212]),
.io_dataIn_213(dataIn[213]),
.io_dataIn_214(dataIn[214]),
.io_dataIn_215(dataIn[215]),
.io_dataIn_216(dataIn[216]),
.io_dataIn_217(dataIn[217]),
.io_dataIn_218(dataIn[218]),
.io_dataIn_219(dataIn[219]),
.io_dataIn_220(dataIn[220]),
.io_dataIn_221(dataIn[221]),
.io_dataIn_222(dataIn[222]),
.io_dataIn_223(dataIn[223]),
.io_dataIn_224(dataIn[224]),
.io_dataIn_225(dataIn[225]),
.io_dataIn_226(dataIn[226]),
.io_dataIn_227(dataIn[227]),
.io_dataIn_228(dataIn[228]),
.io_dataIn_229(dataIn[229]),
.io_dataIn_230(dataIn[230]),
.io_dataIn_231(dataIn[231]),
.io_dataIn_232(dataIn[232]),
.io_dataIn_233(dataIn[233]),
.io_dataIn_234(dataIn[234]),
.io_dataIn_235(dataIn[235]),
.io_dataIn_236(dataIn[236]),
.io_dataIn_237(dataIn[237]),
.io_dataIn_238(dataIn[238]),
.io_dataIn_239(dataIn[239]),
.io_dataIn_240(dataIn[240]),
.io_dataIn_241(dataIn[241]),
.io_dataIn_242(dataIn[242]),
.io_dataIn_243(dataIn[243]),
.io_dataIn_244(dataIn[244]),
.io_dataIn_245(dataIn[245]),
.io_dataIn_246(dataIn[246]),
.io_dataIn_247(dataIn[247]),
.io_dataIn_248(dataIn[248]),
.io_dataIn_249(dataIn[249]),
.io_dataIn_250(dataIn[250]),
.io_dataIn_251(dataIn[251]),
.io_dataIn_252(dataIn[252]),
.io_dataIn_253(dataIn[253]),
.io_dataIn_254(dataIn[254]),
.io_dataIn_255(dataIn[255]),
.io_dataIn_256(dataIn[256]),
.io_dataIn_257(dataIn[257]),
.io_dataIn_258(dataIn[258]),
.io_dataIn_259(dataIn[259]),
.io_dataIn_260(dataIn[260]),
.io_dataIn_261(dataIn[261]),
.io_dataIn_262(dataIn[262]),
.io_dataIn_263(dataIn[263]),
.io_dataIn_264(dataIn[264]),
.io_dataIn_265(dataIn[265]),
.io_dataIn_266(dataIn[266]),
.io_dataIn_267(dataIn[267]),
.io_dataIn_268(dataIn[268]),
.io_dataIn_269(dataIn[269]),
.io_dataIn_270(dataIn[270]),
.io_dataIn_271(dataIn[271]),
.io_dataIn_272(dataIn[272]),
.io_dataIn_273(dataIn[273]),
.io_dataIn_274(dataIn[274]),
.io_dataIn_275(dataIn[275]),
.io_dataIn_276(dataIn[276]),
.io_dataIn_277(dataIn[277]),
.io_dataIn_278(dataIn[278]),
.io_dataIn_279(dataIn[279]),
.io_dataIn_280(dataIn[280]),
.io_dataIn_281(dataIn[281]),
.io_dataIn_282(dataIn[282]),
.io_dataIn_283(dataIn[283]),
.io_dataIn_284(dataIn[284]),
.io_dataIn_285(dataIn[285]),
.io_dataIn_286(dataIn[286]),
.io_dataIn_287(dataIn[287]),
.io_dataIn_288(dataIn[288]),
.io_dataIn_289(dataIn[289]),
.io_dataIn_290(dataIn[290]),
.io_dataIn_291(dataIn[291]),
.io_dataIn_292(dataIn[292]),
.io_dataIn_293(dataIn[293]),
.io_dataIn_294(dataIn[294]),
.io_dataIn_295(dataIn[295]),
.io_dataIn_296(dataIn[296]),
.io_dataIn_297(dataIn[297]),
.io_dataIn_298(dataIn[298]),
.io_dataIn_299(dataIn[299]),
.io_dataIn_300(dataIn[300]),
.io_dataIn_301(dataIn[301]),
.io_dataIn_302(dataIn[302]),
.io_dataIn_303(dataIn[303]),
.io_dataIn_304(dataIn[304]),
.io_dataIn_305(dataIn[305]),
.io_dataIn_306(dataIn[306]),
.io_dataIn_307(dataIn[307]),
.io_dataIn_308(dataIn[308]),
.io_dataIn_309(dataIn[309]),
.io_dataIn_310(dataIn[310]),
.io_dataIn_311(dataIn[311]),
.io_dataIn_312(dataIn[312]),
.io_dataIn_313(dataIn[313]),
.io_dataIn_314(dataIn[314]),
.io_dataIn_315(dataIn[315]),
.io_dataIn_316(dataIn[316]),
.io_dataIn_317(dataIn[317]),
.io_dataIn_318(dataIn[318]),
.io_dataIn_319(dataIn[319]),
.io_dataIn_320(dataIn[320]),
.io_dataIn_321(dataIn[321]),
.io_dataIn_322(dataIn[322]),
.io_dataIn_323(dataIn[323]),
.io_dataIn_324(dataIn[324]),
.io_dataIn_325(dataIn[325]),
.io_dataIn_326(dataIn[326]),
.io_dataIn_327(dataIn[327]),
.io_dataIn_328(dataIn[328]),
.io_dataIn_329(dataIn[329]),
.io_dataIn_330(dataIn[330]),
.io_dataIn_331(dataIn[331]),
.io_dataIn_332(dataIn[332]),
.io_dataIn_333(dataIn[333]),
.io_dataIn_334(dataIn[334]),
.io_dataIn_335(dataIn[335]),
.io_dataIn_336(dataIn[336]),
.io_dataIn_337(dataIn[337]),
.io_dataIn_338(dataIn[338]),
.io_dataIn_339(dataIn[339]),
.io_dataIn_340(dataIn[340]),
.io_dataIn_341(dataIn[341]),
.io_dataIn_342(dataIn[342]),
.io_dataIn_343(dataIn[343]),
.io_dataIn_344(dataIn[344]),
.io_dataIn_345(dataIn[345]),
.io_dataIn_346(dataIn[346]),
.io_dataIn_347(dataIn[347]),
.io_dataIn_348(dataIn[348]),
.io_dataIn_349(dataIn[349]),
.io_dataIn_350(dataIn[350]),
.io_dataIn_351(dataIn[351]),
.io_dataIn_352(dataIn[352]),
.io_dataIn_353(dataIn[353]),
.io_dataIn_354(dataIn[354]),
.io_dataIn_355(dataIn[355]),
.io_dataIn_356(dataIn[356]),
.io_dataIn_357(dataIn[357]),
.io_dataIn_358(dataIn[358]),
.io_dataIn_359(dataIn[359]),
.io_dataIn_360(dataIn[360]),
.io_dataIn_361(dataIn[361]),
.io_dataIn_362(dataIn[362]),
.io_dataIn_363(dataIn[363]),
.io_dataIn_364(dataIn[364]),
.io_dataIn_365(dataIn[365]),
.io_dataIn_366(dataIn[366]),
.io_dataIn_367(dataIn[367]),
.io_dataIn_368(dataIn[368]),
.io_dataIn_369(dataIn[369]),
.io_dataIn_370(dataIn[370]),
.io_dataIn_371(dataIn[371]),
.io_dataIn_372(dataIn[372]),
.io_dataIn_373(dataIn[373]),
.io_dataIn_374(dataIn[374]),
.io_dataIn_375(dataIn[375]),
.io_dataIn_376(dataIn[376]),
.io_dataIn_377(dataIn[377]),
.io_dataIn_378(dataIn[378]),
.io_dataIn_379(dataIn[379]),
.io_dataIn_380(dataIn[380]),
.io_dataIn_381(dataIn[381]),
.io_dataIn_382(dataIn[382]),
.io_dataIn_383(dataIn[383]),
.io_dataIn_384(dataIn[384]),
.io_dataIn_385(dataIn[385]),
.io_dataIn_386(dataIn[386]),
.io_dataIn_387(dataIn[387]),
.io_dataIn_388(dataIn[388]),
.io_dataIn_389(dataIn[389]),
.io_dataIn_390(dataIn[390]),
.io_dataIn_391(dataIn[391]),
.io_dataIn_392(dataIn[392]),
.io_dataIn_393(dataIn[393]),
.io_dataIn_394(dataIn[394]),
.io_dataIn_395(dataIn[395]),
.io_dataIn_396(dataIn[396]),
.io_dataIn_397(dataIn[397]),
.io_dataIn_398(dataIn[398]),
.io_dataIn_399(dataIn[399]),
.io_dataIn_400(dataIn[400]),
.io_dataIn_401(dataIn[401]),
.io_dataIn_402(dataIn[402]),
.io_dataIn_403(dataIn[403]),
.io_dataIn_404(dataIn[404]),
.io_dataIn_405(dataIn[405]),
.io_dataIn_406(dataIn[406]),
.io_dataIn_407(dataIn[407]),
.io_dataIn_408(dataIn[408]),
.io_dataIn_409(dataIn[409]),
.io_dataIn_410(dataIn[410]),
.io_dataIn_411(dataIn[411]),
.io_dataIn_412(dataIn[412]),
.io_dataIn_413(dataIn[413]),
.io_dataIn_414(dataIn[414]),
.io_dataIn_415(dataIn[415]),
.io_dataIn_416(dataIn[416]),
.io_dataIn_417(dataIn[417]),
.io_dataIn_418(dataIn[418]),
.io_dataIn_419(dataIn[419]),
.io_dataIn_420(dataIn[420]),
.io_dataIn_421(dataIn[421]),
.io_dataIn_422(dataIn[422]),
.io_dataIn_423(dataIn[423]),
.io_dataIn_424(dataIn[424]),
.io_dataIn_425(dataIn[425]),
.io_dataIn_426(dataIn[426]),
.io_dataIn_427(dataIn[427]),
.io_dataIn_428(dataIn[428]),
.io_dataIn_429(dataIn[429]),
.io_dataIn_430(dataIn[430]),
.io_dataIn_431(dataIn[431]),
.io_dataIn_432(dataIn[432]),
.io_dataIn_433(dataIn[433]),
.io_dataIn_434(dataIn[434]),
.io_dataIn_435(dataIn[435]),
.io_dataIn_436(dataIn[436]),
.io_dataIn_437(dataIn[437]),
.io_dataIn_438(dataIn[438]),
.io_dataIn_439(dataIn[439]),
.io_dataIn_440(dataIn[440]),
.io_dataIn_441(dataIn[441]),
.io_dataIn_442(dataIn[442]),
.io_dataIn_443(dataIn[443]),
.io_dataIn_444(dataIn[444]),
.io_dataIn_445(dataIn[445]),
.io_dataIn_446(dataIn[446]),
.io_dataIn_447(dataIn[447]),
.io_dataIn_448(dataIn[448]),
.io_dataIn_449(dataIn[449]),
.io_dataIn_450(dataIn[450]),
.io_dataIn_451(dataIn[451]),
.io_dataIn_452(dataIn[452]),
.io_dataIn_453(dataIn[453]),
.io_dataIn_454(dataIn[454]),
.io_dataIn_455(dataIn[455]),
.io_dataIn_456(dataIn[456]),
.io_dataIn_457(dataIn[457]),
.io_dataIn_458(dataIn[458]),
.io_dataIn_459(dataIn[459]),
.io_dataIn_460(dataIn[460]),
.io_dataIn_461(dataIn[461]),
.io_dataIn_462(dataIn[462]),
.io_dataIn_463(dataIn[463]),
.io_dataIn_464(dataIn[464]),
.io_dataIn_465(dataIn[465]),
.io_dataIn_466(dataIn[466]),
.io_dataIn_467(dataIn[467]),
.io_dataIn_468(dataIn[468]),
.io_dataIn_469(dataIn[469]),
.io_dataIn_470(dataIn[470]),
.io_dataIn_471(dataIn[471]),
.io_dataIn_472(dataIn[472]),
.io_dataIn_473(dataIn[473]),
.io_dataIn_474(dataIn[474]),
.io_dataIn_475(dataIn[475]),
.io_dataIn_476(dataIn[476]),
.io_dataIn_477(dataIn[477]),
.io_dataIn_478(dataIn[478]),
.io_dataIn_479(dataIn[479]),
.io_dataIn_480(dataIn[480]),
.io_dataIn_481(dataIn[481]),
.io_dataIn_482(dataIn[482]),
.io_dataIn_483(dataIn[483]),
.io_dataIn_484(dataIn[484]),
.io_dataIn_485(dataIn[485]),
.io_dataIn_486(dataIn[486]),
.io_dataIn_487(dataIn[487]),
.io_dataIn_488(dataIn[488]),
.io_dataIn_489(dataIn[489]),
.io_dataIn_490(dataIn[490]),
.io_dataIn_491(dataIn[491]),
.io_dataIn_492(dataIn[492]),
.io_dataIn_493(dataIn[493]),
.io_dataIn_494(dataIn[494]),
.io_dataIn_495(dataIn[495]),
.io_dataIn_496(dataIn[496]),
.io_dataIn_497(dataIn[497]),
.io_dataIn_498(dataIn[498]),
.io_dataIn_499(dataIn[499]),
.io_dataIn_500(dataIn[500]),
.io_dataIn_501(dataIn[501]),
.io_dataIn_502(dataIn[502]),
.io_dataIn_503(dataIn[503]),
.io_dataIn_504(dataIn[504]),
.io_dataIn_505(dataIn[505]),
.io_dataIn_506(dataIn[506]),
.io_dataIn_507(dataIn[507]),
.io_dataIn_508(dataIn[508]),
.io_dataIn_509(dataIn[509]),
.io_dataIn_510(dataIn[510]),
.io_dataIn_511(dataIn[511]),
.io_dataIn_512(dataIn[512]),
.io_dataIn_513(dataIn[513]),
.io_dataIn_514(dataIn[514]),
.io_dataIn_515(dataIn[515]),
.io_dataIn_516(dataIn[516]),
.io_dataIn_517(dataIn[517]),
.io_dataIn_518(dataIn[518]),
.io_dataIn_519(dataIn[519]),
.io_dataIn_520(dataIn[520]),
.io_dataIn_521(dataIn[521]),
.io_dataIn_522(dataIn[522]),
.io_dataIn_523(dataIn[523]),
.io_dataIn_524(dataIn[524]),
.io_dataIn_525(dataIn[525]),
.io_dataIn_526(dataIn[526]),
.io_dataIn_527(dataIn[527]),
.io_dataIn_528(dataIn[528]),
.io_dataIn_529(dataIn[529]),
.io_dataIn_530(dataIn[530]),
.io_dataIn_531(dataIn[531]),
.io_dataIn_532(dataIn[532]),
.io_dataIn_533(dataIn[533]),
.io_dataIn_534(dataIn[534]),
.io_dataIn_535(dataIn[535]),
.io_dataIn_536(dataIn[536]),
.io_dataIn_537(dataIn[537]),
.io_dataIn_538(dataIn[538]),
.io_dataIn_539(dataIn[539]),
.io_dataIn_540(dataIn[540]),
.io_dataIn_541(dataIn[541]),
.io_dataIn_542(dataIn[542]),
.io_dataIn_543(dataIn[543]),
.io_dataIn_544(dataIn[544]),
.io_dataIn_545(dataIn[545]),
.io_dataIn_546(dataIn[546]),
.io_dataIn_547(dataIn[547]),
.io_dataIn_548(dataIn[548]),
.io_dataIn_549(dataIn[549]),
.io_dataIn_550(dataIn[550]),
.io_dataIn_551(dataIn[551]),
.io_dataIn_552(dataIn[552]),
.io_dataIn_553(dataIn[553]),
.io_dataIn_554(dataIn[554]),
.io_dataIn_555(dataIn[555]),
.io_dataIn_556(dataIn[556]),
.io_dataIn_557(dataIn[557]),
.io_dataIn_558(dataIn[558]),
.io_dataIn_559(dataIn[559]),
.io_dataIn_560(dataIn[560]),
.io_dataIn_561(dataIn[561]),
.io_dataIn_562(dataIn[562]),
.io_dataIn_563(dataIn[563]),
.io_dataIn_564(dataIn[564]),
.io_dataIn_565(dataIn[565]),
.io_dataIn_566(dataIn[566]),
.io_dataIn_567(dataIn[567]),
.io_dataIn_568(dataIn[568]),
.io_dataIn_569(dataIn[569]),
.io_dataIn_570(dataIn[570]),
.io_dataIn_571(dataIn[571]),
.io_dataIn_572(dataIn[572]),
.io_dataIn_573(dataIn[573]),
.io_dataIn_574(dataIn[574]),
.io_dataIn_575(dataIn[575]),
.io_dataIn_576(dataIn[576]),
.io_dataIn_577(dataIn[577]),
.io_dataIn_578(dataIn[578]),
.io_dataIn_579(dataIn[579]),
.io_dataIn_580(dataIn[580]),
.io_dataIn_581(dataIn[581]),
.io_dataIn_582(dataIn[582]),
.io_dataIn_583(dataIn[583]),
.io_dataIn_584(dataIn[584]),
.io_dataIn_585(dataIn[585]),
.io_dataIn_586(dataIn[586]),
.io_dataIn_587(dataIn[587]),
.io_dataIn_588(dataIn[588]),
.io_dataIn_589(dataIn[589]),
.io_dataIn_590(dataIn[590]),
.io_dataIn_591(dataIn[591]),
.io_dataIn_592(dataIn[592]),
.io_dataIn_593(dataIn[593]),
.io_dataIn_594(dataIn[594]),
.io_dataIn_595(dataIn[595]),
.io_dataIn_596(dataIn[596]),
.io_dataIn_597(dataIn[597]),
.io_dataIn_598(dataIn[598]),
.io_dataIn_599(dataIn[599]),
.io_dataIn_600(dataIn[600]),
.io_dataIn_601(dataIn[601]),
.io_dataIn_602(dataIn[602]),
.io_dataIn_603(dataIn[603]),
.io_dataIn_604(dataIn[604]),
.io_dataIn_605(dataIn[605]),
.io_dataIn_606(dataIn[606]),
.io_dataIn_607(dataIn[607]),
.io_dataIn_608(dataIn[608]),
.io_dataIn_609(dataIn[609]),
.io_dataIn_610(dataIn[610]),
.io_dataIn_611(dataIn[611]),
.io_dataIn_612(dataIn[612]),
.io_dataIn_613(dataIn[613]),
.io_dataIn_614(dataIn[614]),
.io_dataIn_615(dataIn[615]),
.io_dataIn_616(dataIn[616]),
.io_dataIn_617(dataIn[617]),
.io_dataIn_618(dataIn[618]),
.io_dataIn_619(dataIn[619]),
.io_dataIn_620(dataIn[620]),
.io_dataIn_621(dataIn[621]),
.io_dataIn_622(dataIn[622]),
.io_dataIn_623(dataIn[623]),
.io_dataIn_624(dataIn[624]),
.io_dataIn_625(dataIn[625]),
.io_dataIn_626(dataIn[626]),
.io_dataIn_627(dataIn[627]),
.io_dataIn_628(dataIn[628]),
.io_dataIn_629(dataIn[629]),
.io_dataIn_630(dataIn[630]),
.io_dataIn_631(dataIn[631]),
.io_dataIn_632(dataIn[632]),
.io_dataIn_633(dataIn[633]),
.io_dataIn_634(dataIn[634]),
.io_dataIn_635(dataIn[635]),
.io_dataIn_636(dataIn[636]),
.io_dataIn_637(dataIn[637]),
.io_dataIn_638(dataIn[638]),
.io_dataIn_639(dataIn[639]),
.io_dataIn_640(dataIn[640]),
.io_dataIn_641(dataIn[641]),
.io_dataIn_642(dataIn[642]),
.io_dataIn_643(dataIn[643]),
.io_dataIn_644(dataIn[644]),
.io_dataIn_645(dataIn[645]),
.io_dataIn_646(dataIn[646]),
.io_dataIn_647(dataIn[647]),
.io_dataIn_648(dataIn[648]),
.io_dataIn_649(dataIn[649]),
.io_dataIn_650(dataIn[650]),
.io_dataIn_651(dataIn[651]),
.io_dataIn_652(dataIn[652]),
.io_dataIn_653(dataIn[653]),
.io_dataIn_654(dataIn[654]),
.io_dataIn_655(dataIn[655]),
.io_dataIn_656(dataIn[656]),
.io_dataIn_657(dataIn[657]),
.io_dataIn_658(dataIn[658]),
.io_dataIn_659(dataIn[659]),
.io_dataIn_660(dataIn[660]),
.io_dataIn_661(dataIn[661]),
.io_dataIn_662(dataIn[662]),
.io_dataIn_663(dataIn[663]),
.io_dataIn_664(dataIn[664]),
.io_dataIn_665(dataIn[665]),
.io_dataIn_666(dataIn[666]),
.io_dataIn_667(dataIn[667]),
.io_dataIn_668(dataIn[668]),
.io_dataIn_669(dataIn[669]),
.io_dataIn_670(dataIn[670]),
.io_dataIn_671(dataIn[671]),
.io_dataIn_672(dataIn[672]),
.io_dataIn_673(dataIn[673]),
.io_dataIn_674(dataIn[674]),
.io_dataIn_675(dataIn[675]),
.io_dataIn_676(dataIn[676]),
.io_dataIn_677(dataIn[677]),
.io_dataIn_678(dataIn[678]),
.io_dataIn_679(dataIn[679]),
.io_dataIn_680(dataIn[680]),
.io_dataIn_681(dataIn[681]),
.io_dataIn_682(dataIn[682]),
.io_dataIn_683(dataIn[683]),
.io_dataIn_684(dataIn[684]),
.io_dataIn_685(dataIn[685]),
.io_dataIn_686(dataIn[686]),
.io_dataIn_687(dataIn[687]),
.io_dataIn_688(dataIn[688]),
.io_dataIn_689(dataIn[689]),
.io_dataIn_690(dataIn[690]),
.io_dataIn_691(dataIn[691]),
.io_dataIn_692(dataIn[692]),
.io_dataIn_693(dataIn[693]),
.io_dataIn_694(dataIn[694]),
.io_dataIn_695(dataIn[695]),
.io_dataIn_696(dataIn[696]),
.io_dataIn_697(dataIn[697]),
.io_dataIn_698(dataIn[698]),
.io_dataIn_699(dataIn[699]),
.io_dataIn_700(dataIn[700]),
.io_dataIn_701(dataIn[701]),
.io_dataIn_702(dataIn[702]),
.io_dataIn_703(dataIn[703]),
.io_dataIn_704(dataIn[704]),
.io_dataIn_705(dataIn[705]),
.io_dataIn_706(dataIn[706]),
.io_dataIn_707(dataIn[707]),
.io_dataIn_708(dataIn[708]),
.io_dataIn_709(dataIn[709]),
.io_dataIn_710(dataIn[710]),
.io_dataIn_711(dataIn[711]),
.io_dataIn_712(dataIn[712]),
.io_dataIn_713(dataIn[713]),
.io_dataIn_714(dataIn[714]),
.io_dataIn_715(dataIn[715]),
.io_dataIn_716(dataIn[716]),
.io_dataIn_717(dataIn[717]),
.io_dataIn_718(dataIn[718]),
.io_dataIn_719(dataIn[719]),
.io_dataIn_720(dataIn[720]),
.io_dataIn_721(dataIn[721]),
.io_dataIn_722(dataIn[722]),
.io_dataIn_723(dataIn[723]),
.io_dataIn_724(dataIn[724]),
.io_dataIn_725(dataIn[725]),
.io_dataIn_726(dataIn[726]),
.io_dataIn_727(dataIn[727]),
.io_dataIn_728(dataIn[728]),
.io_dataIn_729(dataIn[729]),
.io_dataIn_730(dataIn[730]),
.io_dataIn_731(dataIn[731]),
.io_dataIn_732(dataIn[732]),
.io_dataIn_733(dataIn[733]),
.io_dataIn_734(dataIn[734]),
.io_dataIn_735(dataIn[735]),
.io_dataIn_736(dataIn[736]),
.io_dataIn_737(dataIn[737]),
.io_dataIn_738(dataIn[738]),
.io_dataIn_739(dataIn[739]),
.io_dataIn_740(dataIn[740]),
.io_dataIn_741(dataIn[741]),
.io_dataIn_742(dataIn[742]),
.io_dataIn_743(dataIn[743]),
.io_dataIn_744(dataIn[744]),
.io_dataIn_745(dataIn[745]),
.io_dataIn_746(dataIn[746]),
.io_dataIn_747(dataIn[747]),
.io_dataIn_748(dataIn[748]),
.io_dataIn_749(dataIn[749]),
.io_dataIn_750(dataIn[750]),
.io_dataIn_751(dataIn[751]),
.io_dataIn_752(dataIn[752]),
.io_dataIn_753(dataIn[753]),
.io_dataIn_754(dataIn[754]),
.io_dataIn_755(dataIn[755]),
.io_dataIn_756(dataIn[756]),
.io_dataIn_757(dataIn[757]),
.io_dataIn_758(dataIn[758]),
.io_dataIn_759(dataIn[759]),
.io_dataIn_760(dataIn[760]),
.io_dataIn_761(dataIn[761]),
.io_dataIn_762(dataIn[762]),
.io_dataIn_763(dataIn[763]),
.io_dataIn_764(dataIn[764]),
.io_dataIn_765(dataIn[765]),
.io_dataIn_766(dataIn[766]),
.io_dataIn_767(dataIn[767]),
.io_dataIn_768(dataIn[768]),
.io_dataIn_769(dataIn[769]),
.io_dataIn_770(dataIn[770]),
.io_dataIn_771(dataIn[771]),
.io_dataIn_772(dataIn[772]),
.io_dataIn_773(dataIn[773]),
.io_dataIn_774(dataIn[774]),
.io_dataIn_775(dataIn[775]),
.io_dataIn_776(dataIn[776]),
.io_dataIn_777(dataIn[777]),
.io_dataIn_778(dataIn[778]),
.io_dataIn_779(dataIn[779]),
.io_dataIn_780(dataIn[780]),
.io_dataIn_781(dataIn[781]),
.io_dataIn_782(dataIn[782]),
.io_dataIn_783(dataIn[783]),
.io_dataIn_784(dataIn[784]),
.io_dataIn_785(dataIn[785]),
.io_dataIn_786(dataIn[786]),
.io_dataIn_787(dataIn[787]),
.io_dataIn_788(dataIn[788]),
.io_dataIn_789(dataIn[789]),
.io_dataIn_790(dataIn[790]),
.io_dataIn_791(dataIn[791]),
.io_dataIn_792(dataIn[792]),
.io_dataIn_793(dataIn[793]),
.io_dataIn_794(dataIn[794]),
.io_dataIn_795(dataIn[795]),
.io_dataIn_796(dataIn[796]),
.io_dataIn_797(dataIn[797]),
.io_dataIn_798(dataIn[798]),
.io_dataIn_799(dataIn[799]),
.io_dataIn_800(dataIn[800]),
.io_dataIn_801(dataIn[801]),
.io_dataIn_802(dataIn[802]),
.io_dataIn_803(dataIn[803]),
.io_dataIn_804(dataIn[804]),
.io_dataIn_805(dataIn[805]),
.io_dataIn_806(dataIn[806]),
.io_dataIn_807(dataIn[807]),
.io_dataIn_808(dataIn[808]),
.io_dataIn_809(dataIn[809]),
.io_dataIn_810(dataIn[810]),
.io_dataIn_811(dataIn[811]),
.io_dataIn_812(dataIn[812]),
.io_dataIn_813(dataIn[813]),
.io_dataIn_814(dataIn[814]),
.io_dataIn_815(dataIn[815]),
.io_dataIn_816(dataIn[816]),
.io_dataIn_817(dataIn[817]),
.io_dataIn_818(dataIn[818]),
.io_dataIn_819(dataIn[819]),
.io_dataIn_820(dataIn[820]),
.io_dataIn_821(dataIn[821]),
.io_dataIn_822(dataIn[822]),
.io_dataIn_823(dataIn[823]),
.io_dataIn_824(dataIn[824]),
.io_dataIn_825(dataIn[825]),
.io_dataIn_826(dataIn[826]),
.io_dataIn_827(dataIn[827]),
.io_dataIn_828(dataIn[828]),
.io_dataIn_829(dataIn[829]),
.io_dataIn_830(dataIn[830]),
.io_dataIn_831(dataIn[831]),
.io_dataIn_832(dataIn[832]),
.io_dataIn_833(dataIn[833]),
.io_dataIn_834(dataIn[834]),
.io_dataIn_835(dataIn[835]),
.io_dataIn_836(dataIn[836]),
.io_dataIn_837(dataIn[837]),
.io_dataIn_838(dataIn[838]),
.io_dataIn_839(dataIn[839]),
.io_dataIn_840(dataIn[840]),
.io_dataIn_841(dataIn[841]),
.io_dataIn_842(dataIn[842]),
.io_dataIn_843(dataIn[843]),
.io_dataIn_844(dataIn[844]),
.io_dataIn_845(dataIn[845]),
.io_dataIn_846(dataIn[846]),
.io_dataIn_847(dataIn[847]),
.io_dataIn_848(dataIn[848]),
.io_dataIn_849(dataIn[849]),
.io_dataIn_850(dataIn[850]),
.io_dataIn_851(dataIn[851]),
.io_dataIn_852(dataIn[852]),
.io_dataIn_853(dataIn[853]),
.io_dataIn_854(dataIn[854]),
.io_dataIn_855(dataIn[855]),
.io_dataIn_856(dataIn[856]),
.io_dataIn_857(dataIn[857]),
.io_dataIn_858(dataIn[858]),
.io_dataIn_859(dataIn[859]),
.io_dataIn_860(dataIn[860]),
.io_dataIn_861(dataIn[861]),
.io_dataIn_862(dataIn[862]),
.io_dataIn_863(dataIn[863]),
.io_dataIn_864(dataIn[864]),
.io_dataIn_865(dataIn[865]),
.io_dataIn_866(dataIn[866]),
.io_dataIn_867(dataIn[867]),
.io_dataIn_868(dataIn[868]),
.io_dataIn_869(dataIn[869]),
.io_dataIn_870(dataIn[870]),
.io_dataIn_871(dataIn[871]),
.io_dataIn_872(dataIn[872]),
.io_dataIn_873(dataIn[873]),
.io_dataIn_874(dataIn[874]),
.io_dataIn_875(dataIn[875]),
.io_dataIn_876(dataIn[876]),
.io_dataIn_877(dataIn[877]),
.io_dataIn_878(dataIn[878]),
.io_dataIn_879(dataIn[879]),
.io_dataIn_880(dataIn[880]),
.io_dataIn_881(dataIn[881]),
.io_dataIn_882(dataIn[882]),
.io_dataIn_883(dataIn[883]),
.io_dataIn_884(dataIn[884]),
.io_dataIn_885(dataIn[885]),
.io_dataIn_886(dataIn[886]),
.io_dataIn_887(dataIn[887]),
.io_dataIn_888(dataIn[888]),
.io_dataIn_889(dataIn[889]),
.io_dataIn_890(dataIn[890]),
.io_dataIn_891(dataIn[891]),
.io_dataIn_892(dataIn[892]),
.io_dataIn_893(dataIn[893]),
.io_dataIn_894(dataIn[894]),
.io_dataIn_895(dataIn[895]),
.io_dataIn_896(dataIn[896]),
.io_dataIn_897(dataIn[897]),
.io_dataIn_898(dataIn[898]),
.io_dataIn_899(dataIn[899]),
.io_dataIn_900(dataIn[900]),
.io_dataIn_901(dataIn[901]),
.io_dataIn_902(dataIn[902]),
.io_dataIn_903(dataIn[903]),
.io_dataIn_904(dataIn[904]),
.io_dataIn_905(dataIn[905]),
.io_dataIn_906(dataIn[906]),
.io_dataIn_907(dataIn[907]),
.io_dataIn_908(dataIn[908]),
.io_dataIn_909(dataIn[909]),
.io_dataIn_910(dataIn[910]),
.io_dataIn_911(dataIn[911]),
.io_dataIn_912(dataIn[912]),
.io_dataIn_913(dataIn[913]),
.io_dataIn_914(dataIn[914]),
.io_dataIn_915(dataIn[915]),
.io_dataIn_916(dataIn[916]),
.io_dataIn_917(dataIn[917]),
.io_dataIn_918(dataIn[918]),
.io_dataIn_919(dataIn[919]),
.io_dataIn_920(dataIn[920]),
.io_dataIn_921(dataIn[921]),
.io_dataIn_922(dataIn[922]),
.io_dataIn_923(dataIn[923]),
.io_dataIn_924(dataIn[924]),
.io_dataIn_925(dataIn[925]),
.io_dataIn_926(dataIn[926]),
.io_dataIn_927(dataIn[927]),
.io_dataIn_928(dataIn[928]),
.io_dataIn_929(dataIn[929]),
.io_dataIn_930(dataIn[930]),
.io_dataIn_931(dataIn[931]),
.io_dataIn_932(dataIn[932]),
.io_dataIn_933(dataIn[933]),
.io_dataIn_934(dataIn[934]),
.io_dataIn_935(dataIn[935]),
.io_dataIn_936(dataIn[936]),
.io_dataIn_937(dataIn[937]),
.io_dataIn_938(dataIn[938]),
.io_dataIn_939(dataIn[939]),
.io_dataIn_940(dataIn[940]),
.io_dataIn_941(dataIn[941]),
.io_dataIn_942(dataIn[942]),
.io_dataIn_943(dataIn[943]),
.io_dataIn_944(dataIn[944]),
.io_dataIn_945(dataIn[945]),
.io_dataIn_946(dataIn[946]),
.io_dataIn_947(dataIn[947]),
.io_dataIn_948(dataIn[948]),
.io_dataIn_949(dataIn[949]),
.io_dataIn_950(dataIn[950]),
.io_dataIn_951(dataIn[951]),
.io_dataIn_952(dataIn[952]),
.io_dataIn_953(dataIn[953]),
.io_dataIn_954(dataIn[954]),
.io_dataIn_955(dataIn[955]),
.io_dataIn_956(dataIn[956]),
.io_dataIn_957(dataIn[957]),
.io_dataIn_958(dataIn[958]),
.io_dataIn_959(dataIn[959]),
.io_dataIn_960(dataIn[960]),
.io_dataIn_961(dataIn[961]),
.io_dataIn_962(dataIn[962]),
.io_dataIn_963(dataIn[963]),
.io_dataIn_964(dataIn[964]),
.io_dataIn_965(dataIn[965]),
.io_dataIn_966(dataIn[966]),
.io_dataIn_967(dataIn[967]),
.io_dataIn_968(dataIn[968]),
.io_dataIn_969(dataIn[969]),
.io_dataIn_970(dataIn[970]),
.io_dataIn_971(dataIn[971]),
.io_dataIn_972(dataIn[972]),
.io_dataIn_973(dataIn[973]),
.io_dataIn_974(dataIn[974]),
.io_dataIn_975(dataIn[975]),
.io_dataIn_976(dataIn[976]),
.io_dataIn_977(dataIn[977]),
.io_dataIn_978(dataIn[978]),
.io_dataIn_979(dataIn[979]),
.io_dataIn_980(dataIn[980]),
.io_dataIn_981(dataIn[981]),
.io_dataIn_982(dataIn[982]),
.io_dataIn_983(dataIn[983]),
.io_dataIn_984(dataIn[984]),
.io_dataIn_985(dataIn[985]),
.io_dataIn_986(dataIn[986]),
.io_dataIn_987(dataIn[987]),
.io_dataIn_988(dataIn[988]),
.io_dataIn_989(dataIn[989]),
.io_dataIn_990(dataIn[990]),
.io_dataIn_991(dataIn[991]),
.io_dataIn_992(dataIn[992]),
.io_dataIn_993(dataIn[993]),
.io_dataIn_994(dataIn[994]),
.io_dataIn_995(dataIn[995]),
.io_dataIn_996(dataIn[996]),
.io_dataIn_997(dataIn[997]),
.io_dataIn_998(dataIn[998]),
.io_dataIn_999(dataIn[999]),
.io_dataIn_1000(dataIn[1000]),
.io_dataIn_1001(dataIn[1001]),
.io_dataIn_1002(dataIn[1002]),
.io_dataIn_1003(dataIn[1003]),
.io_dataIn_1004(dataIn[1004]),
.io_dataIn_1005(dataIn[1005]),
.io_dataIn_1006(dataIn[1006]),
.io_dataIn_1007(dataIn[1007]),
.io_dataIn_1008(dataIn[1008]),
.io_dataIn_1009(dataIn[1009]),
.io_dataIn_1010(dataIn[1010]),
.io_dataIn_1011(dataIn[1011]),
.io_dataIn_1012(dataIn[1012]),
.io_dataIn_1013(dataIn[1013]),
.io_dataIn_1014(dataIn[1014]),
.io_dataIn_1015(dataIn[1015]),
.io_dataIn_1016(dataIn[1016]),
.io_dataIn_1017(dataIn[1017]),
.io_dataIn_1018(dataIn[1018]),
.io_dataIn_1019(dataIn[1019]),
.io_dataIn_1020(dataIn[1020]),
.io_dataIn_1021(dataIn[1021]),
.io_dataIn_1022(dataIn[1022]),
.io_dataIn_1023(dataIn[1023]),
.io_dataIn_1024(dataIn[1024]),
.io_dataIn_1025(dataIn[1025]),
.io_dataIn_1026(dataIn[1026]),
.io_dataIn_1027(dataIn[1027]),
.io_dataIn_1028(dataIn[1028]),
.io_dataIn_1029(dataIn[1029]),
.io_dataIn_1030(dataIn[1030]),
.io_dataIn_1031(dataIn[1031]),
.io_dataIn_1032(dataIn[1032]),
.io_dataIn_1033(dataIn[1033]),
.io_dataIn_1034(dataIn[1034]),
.io_dataIn_1035(dataIn[1035]),
.io_dataIn_1036(dataIn[1036]),
.io_dataIn_1037(dataIn[1037]),
.io_dataIn_1038(dataIn[1038]),
.io_dataIn_1039(dataIn[1039]),
.io_dataIn_1040(dataIn[1040]),
.io_dataIn_1041(dataIn[1041]),
.io_dataIn_1042(dataIn[1042]),
.io_dataIn_1043(dataIn[1043]),
.io_dataIn_1044(dataIn[1044]),
.io_dataIn_1045(dataIn[1045]),
.io_dataIn_1046(dataIn[1046]),
.io_dataIn_1047(dataIn[1047]),
.io_dataIn_1048(dataIn[1048]),
.io_dataIn_1049(dataIn[1049]),
.io_dataIn_1050(dataIn[1050]),
.io_dataIn_1051(dataIn[1051]),
.io_dataIn_1052(dataIn[1052]),
.io_dataIn_1053(dataIn[1053]),
.io_dataIn_1054(dataIn[1054]),
.io_dataIn_1055(dataIn[1055]),
.io_dataIn_1056(dataIn[1056]),
.io_dataIn_1057(dataIn[1057]),
.io_dataIn_1058(dataIn[1058]),
.io_dataIn_1059(dataIn[1059]),
.io_dataIn_1060(dataIn[1060]),
.io_dataIn_1061(dataIn[1061]),
.io_dataIn_1062(dataIn[1062]),
.io_dataIn_1063(dataIn[1063]),
.io_dataIn_1064(dataIn[1064]),
.io_dataIn_1065(dataIn[1065]),
.io_dataIn_1066(dataIn[1066]),
.io_dataIn_1067(dataIn[1067]),
.io_dataIn_1068(dataIn[1068]),
.io_dataIn_1069(dataIn[1069]),
.io_dataIn_1070(dataIn[1070]),
.io_dataIn_1071(dataIn[1071]),
.io_dataIn_1072(dataIn[1072]),
.io_dataIn_1073(dataIn[1073]),
.io_dataIn_1074(dataIn[1074]),
.io_dataIn_1075(dataIn[1075]),
.io_dataIn_1076(dataIn[1076]),
.io_dataIn_1077(dataIn[1077]),
.io_dataIn_1078(dataIn[1078]),
.io_dataIn_1079(dataIn[1079]),
.io_dataIn_1080(dataIn[1080]),
.io_dataIn_1081(dataIn[1081]),
.io_dataIn_1082(dataIn[1082]),
.io_dataIn_1083(dataIn[1083]),
.io_dataIn_1084(dataIn[1084]),
.io_dataIn_1085(dataIn[1085]),
.io_dataIn_1086(dataIn[1086]),
.io_dataIn_1087(dataIn[1087]),
.io_dataIn_1088(dataIn[1088]),
.io_dataIn_1089(dataIn[1089]),
.io_dataIn_1090(dataIn[1090]),
.io_dataIn_1091(dataIn[1091]),
.io_dataIn_1092(dataIn[1092]),
.io_dataIn_1093(dataIn[1093]),
.io_dataIn_1094(dataIn[1094]),
.io_dataIn_1095(dataIn[1095]),
.io_dataIn_1096(dataIn[1096]),
.io_dataIn_1097(dataIn[1097]),
.io_dataIn_1098(dataIn[1098]),
.io_dataIn_1099(dataIn[1099]),
.io_dataIn_1100(dataIn[1100]),
.io_dataIn_1101(dataIn[1101]),
.io_dataIn_1102(dataIn[1102]),
.io_dataIn_1103(dataIn[1103]),
.io_dataIn_1104(dataIn[1104]),
.io_dataIn_1105(dataIn[1105]),
.io_dataIn_1106(dataIn[1106]),
.io_dataIn_1107(dataIn[1107]),
.io_dataIn_1108(dataIn[1108]),
.io_dataIn_1109(dataIn[1109]),
.io_dataIn_1110(dataIn[1110]),
.io_dataIn_1111(dataIn[1111]),
.io_dataIn_1112(dataIn[1112]),
.io_dataIn_1113(dataIn[1113]),
.io_dataIn_1114(dataIn[1114]),
.io_dataIn_1115(dataIn[1115]),
.io_dataIn_1116(dataIn[1116]),
.io_dataIn_1117(dataIn[1117]),
.io_dataIn_1118(dataIn[1118]),
.io_dataIn_1119(dataIn[1119]),
.io_dataIn_1120(dataIn[1120]),
.io_dataIn_1121(dataIn[1121]),
.io_dataIn_1122(dataIn[1122]),
.io_dataIn_1123(dataIn[1123]),
.io_dataIn_1124(dataIn[1124]),
.io_dataIn_1125(dataIn[1125]),
.io_dataIn_1126(dataIn[1126]),
.io_dataIn_1127(dataIn[1127]),
.io_dataIn_1128(dataIn[1128]),
.io_dataIn_1129(dataIn[1129]),
.io_dataIn_1130(dataIn[1130]),
.io_dataIn_1131(dataIn[1131]),
.io_dataIn_1132(dataIn[1132]),
.io_dataIn_1133(dataIn[1133]),
.io_dataIn_1134(dataIn[1134]),
.io_dataIn_1135(dataIn[1135]),
.io_dataIn_1136(dataIn[1136]),
.io_dataIn_1137(dataIn[1137]),
.io_dataIn_1138(dataIn[1138]),
.io_dataIn_1139(dataIn[1139]),
.io_dataIn_1140(dataIn[1140]),
.io_dataIn_1141(dataIn[1141]),
.io_dataIn_1142(dataIn[1142]),
.io_dataIn_1143(dataIn[1143]),
.io_dataIn_1144(dataIn[1144]),
.io_dataIn_1145(dataIn[1145]),
.io_dataIn_1146(dataIn[1146]),
.io_dataIn_1147(dataIn[1147]),
.io_dataIn_1148(dataIn[1148]),
.io_dataIn_1149(dataIn[1149]),
.io_dataIn_1150(dataIn[1150]),
.io_dataIn_1151(dataIn[1151]),
.io_dataIn_1152(dataIn[1152]),
.io_dataIn_1153(dataIn[1153]),
.io_dataIn_1154(dataIn[1154]),
.io_dataIn_1155(dataIn[1155]),
.io_dataIn_1156(dataIn[1156]),
.io_dataIn_1157(dataIn[1157]),
.io_dataIn_1158(dataIn[1158]),
.io_dataIn_1159(dataIn[1159]),
.io_dataIn_1160(dataIn[1160]),
.io_dataIn_1161(dataIn[1161]),
.io_dataIn_1162(dataIn[1162]),
.io_dataIn_1163(dataIn[1163]),
.io_dataIn_1164(dataIn[1164]),
.io_dataIn_1165(dataIn[1165]),
.io_dataIn_1166(dataIn[1166]),
.io_dataIn_1167(dataIn[1167]),
.io_dataIn_1168(dataIn[1168]),
.io_dataIn_1169(dataIn[1169]),
.io_dataIn_1170(dataIn[1170]),
.io_dataIn_1171(dataIn[1171]),
.io_dataIn_1172(dataIn[1172]),
.io_dataIn_1173(dataIn[1173]),
.io_dataIn_1174(dataIn[1174]),
.io_dataIn_1175(dataIn[1175]),
.io_dataIn_1176(dataIn[1176]),
.io_dataIn_1177(dataIn[1177]),
.io_dataIn_1178(dataIn[1178]),
.io_dataIn_1179(dataIn[1179]),
.io_dataIn_1180(dataIn[1180]),
.io_dataIn_1181(dataIn[1181]),
.io_dataIn_1182(dataIn[1182]),
.io_dataIn_1183(dataIn[1183]),
.io_dataIn_1184(dataIn[1184]),
.io_dataIn_1185(dataIn[1185]),
.io_dataIn_1186(dataIn[1186]),
.io_dataIn_1187(dataIn[1187]),
.io_dataIn_1188(dataIn[1188]),
.io_dataIn_1189(dataIn[1189]),
.io_dataIn_1190(dataIn[1190]),
.io_dataIn_1191(dataIn[1191]),
.io_dataIn_1192(dataIn[1192]),
.io_dataIn_1193(dataIn[1193]),
.io_dataIn_1194(dataIn[1194]),
.io_dataIn_1195(dataIn[1195]),
.io_dataIn_1196(dataIn[1196]),
.io_dataIn_1197(dataIn[1197]),
.io_dataIn_1198(dataIn[1198]),
.io_dataIn_1199(dataIn[1199]),
.io_dataIn_1200(dataIn[1200]),
.io_dataIn_1201(dataIn[1201]),
.io_dataIn_1202(dataIn[1202]),
.io_dataIn_1203(dataIn[1203]),
.io_dataIn_1204(dataIn[1204]),
.io_dataIn_1205(dataIn[1205]),
.io_dataIn_1206(dataIn[1206]),
.io_dataIn_1207(dataIn[1207]),
.io_dataIn_1208(dataIn[1208]),
.io_dataIn_1209(dataIn[1209]),
.io_dataIn_1210(dataIn[1210]),
.io_dataIn_1211(dataIn[1211]),
.io_dataIn_1212(dataIn[1212]),
.io_dataIn_1213(dataIn[1213]),
.io_dataIn_1214(dataIn[1214]),
.io_dataIn_1215(dataIn[1215]),
.io_dataIn_1216(dataIn[1216]),
.io_dataIn_1217(dataIn[1217]),
.io_dataIn_1218(dataIn[1218]),
.io_dataIn_1219(dataIn[1219]),
.io_dataIn_1220(dataIn[1220]),
.io_dataIn_1221(dataIn[1221]),
.io_dataIn_1222(dataIn[1222]),
.io_dataIn_1223(dataIn[1223]),
.io_dataIn_1224(dataIn[1224]),
.io_dataIn_1225(dataIn[1225]),
.io_dataIn_1226(dataIn[1226]),
.io_dataIn_1227(dataIn[1227]),
.io_dataIn_1228(dataIn[1228]),
.io_dataIn_1229(dataIn[1229]),
.io_dataIn_1230(dataIn[1230]),
.io_dataIn_1231(dataIn[1231]),
.io_dataIn_1232(dataIn[1232]),
.io_dataIn_1233(dataIn[1233]),
.io_dataIn_1234(dataIn[1234]),
.io_dataIn_1235(dataIn[1235]),
.io_dataIn_1236(dataIn[1236]),
.io_dataIn_1237(dataIn[1237]),
.io_dataIn_1238(dataIn[1238]),
.io_dataIn_1239(dataIn[1239]),
.io_dataIn_1240(dataIn[1240]),
.io_dataIn_1241(dataIn[1241]),
.io_dataIn_1242(dataIn[1242]),
.io_dataIn_1243(dataIn[1243]),
.io_dataIn_1244(dataIn[1244]),
.io_dataIn_1245(dataIn[1245]),
.io_dataIn_1246(dataIn[1246]),
.io_dataIn_1247(dataIn[1247]),
.io_dataIn_1248(dataIn[1248]),
.io_dataIn_1249(dataIn[1249]),
.io_dataIn_1250(dataIn[1250]),
.io_dataIn_1251(dataIn[1251]),
.io_dataIn_1252(dataIn[1252]),
.io_dataIn_1253(dataIn[1253]),
.io_dataIn_1254(dataIn[1254]),
.io_dataIn_1255(dataIn[1255]),
.io_dataIn_1256(dataIn[1256]),
.io_dataIn_1257(dataIn[1257]),
.io_dataIn_1258(dataIn[1258]),
.io_dataIn_1259(dataIn[1259]),
.io_dataIn_1260(dataIn[1260]),
.io_dataIn_1261(dataIn[1261]),
.io_dataIn_1262(dataIn[1262]),
.io_dataIn_1263(dataIn[1263]),
.io_dataIn_1264(dataIn[1264]),
.io_dataIn_1265(dataIn[1265]),
.io_dataIn_1266(dataIn[1266]),
.io_dataIn_1267(dataIn[1267]),
.io_dataIn_1268(dataIn[1268]),
.io_dataIn_1269(dataIn[1269]),
.io_dataIn_1270(dataIn[1270]),
.io_dataIn_1271(dataIn[1271]),
.io_dataIn_1272(dataIn[1272]),
.io_dataIn_1273(dataIn[1273]),
.io_dataIn_1274(dataIn[1274]),
.io_dataIn_1275(dataIn[1275]),
.io_dataIn_1276(dataIn[1276]),
.io_dataIn_1277(dataIn[1277]),
.io_dataIn_1278(dataIn[1278]),
.io_dataIn_1279(dataIn[1279]),
.io_dataIn_1280(dataIn[1280]),
.io_dataIn_1281(dataIn[1281]),
.io_dataIn_1282(dataIn[1282]),
.io_dataIn_1283(dataIn[1283]),
.io_dataIn_1284(dataIn[1284]),
.io_dataIn_1285(dataIn[1285]),
.io_dataIn_1286(dataIn[1286]),
.io_dataIn_1287(dataIn[1287]),
.io_dataIn_1288(dataIn[1288]),
.io_dataIn_1289(dataIn[1289]),
.io_dataIn_1290(dataIn[1290]),
.io_dataIn_1291(dataIn[1291]),
.io_dataIn_1292(dataIn[1292]),
.io_dataIn_1293(dataIn[1293]),
.io_dataIn_1294(dataIn[1294]),
.io_dataIn_1295(dataIn[1295]),
.io_dataIn_1296(dataIn[1296]),
.io_dataIn_1297(dataIn[1297]),
.io_dataIn_1298(dataIn[1298]),
.io_dataIn_1299(dataIn[1299]),
.io_dataIn_1300(dataIn[1300]),
.io_dataIn_1301(dataIn[1301]),
.io_dataIn_1302(dataIn[1302]),
.io_dataIn_1303(dataIn[1303]),
.io_dataIn_1304(dataIn[1304]),
.io_dataIn_1305(dataIn[1305]),
.io_dataIn_1306(dataIn[1306]),
.io_dataIn_1307(dataIn[1307]),
.io_dataIn_1308(dataIn[1308]),
.io_dataIn_1309(dataIn[1309]),
.io_dataIn_1310(dataIn[1310]),
.io_dataIn_1311(dataIn[1311]),
.io_dataIn_1312(dataIn[1312]),
.io_dataIn_1313(dataIn[1313]),
.io_dataIn_1314(dataIn[1314]),
.io_dataIn_1315(dataIn[1315]),
.io_dataIn_1316(dataIn[1316]),
.io_dataIn_1317(dataIn[1317]),
.io_dataIn_1318(dataIn[1318]),
.io_dataIn_1319(dataIn[1319]),
.io_dataIn_1320(dataIn[1320]),
.io_dataIn_1321(dataIn[1321]),
.io_dataIn_1322(dataIn[1322]),
.io_dataIn_1323(dataIn[1323]),
.io_dataIn_1324(dataIn[1324]),
.io_dataIn_1325(dataIn[1325]),
.io_dataIn_1326(dataIn[1326]),
.io_dataIn_1327(dataIn[1327]),
.io_dataIn_1328(dataIn[1328]),
.io_dataIn_1329(dataIn[1329]),
.io_dataIn_1330(dataIn[1330]),
.io_dataIn_1331(dataIn[1331]),
.io_dataIn_1332(dataIn[1332]),
.io_dataIn_1333(dataIn[1333]),
.io_dataIn_1334(dataIn[1334]),
.io_dataIn_1335(dataIn[1335]),
.io_dataIn_1336(dataIn[1336]),
.io_dataIn_1337(dataIn[1337]),
.io_dataIn_1338(dataIn[1338]),
.io_dataIn_1339(dataIn[1339]),
.io_dataIn_1340(dataIn[1340]),
.io_dataIn_1341(dataIn[1341]),
.io_dataIn_1342(dataIn[1342]),
.io_dataIn_1343(dataIn[1343]),
.io_dataIn_1344(dataIn[1344]),
.io_dataIn_1345(dataIn[1345]),
.io_dataIn_1346(dataIn[1346]),
.io_dataIn_1347(dataIn[1347]),
.io_dataIn_1348(dataIn[1348]),
.io_dataIn_1349(dataIn[1349]),
.io_dataIn_1350(dataIn[1350]),
.io_dataIn_1351(dataIn[1351]),
.io_dataIn_1352(dataIn[1352]),
.io_dataIn_1353(dataIn[1353]),
.io_dataIn_1354(dataIn[1354]),
.io_dataIn_1355(dataIn[1355]),
.io_dataIn_1356(dataIn[1356]),
.io_dataIn_1357(dataIn[1357]),
.io_dataIn_1358(dataIn[1358]),
.io_dataIn_1359(dataIn[1359]),
.io_dataIn_1360(dataIn[1360]),
.io_dataIn_1361(dataIn[1361]),
.io_dataIn_1362(dataIn[1362]),
.io_dataIn_1363(dataIn[1363]),
.io_dataIn_1364(dataIn[1364]),
.io_dataIn_1365(dataIn[1365]),
.io_dataIn_1366(dataIn[1366]),
.io_dataIn_1367(dataIn[1367]),
.io_dataIn_1368(dataIn[1368]),
.io_dataIn_1369(dataIn[1369]),
.io_dataIn_1370(dataIn[1370]),
.io_dataIn_1371(dataIn[1371]),
.io_dataIn_1372(dataIn[1372]),
.io_dataIn_1373(dataIn[1373]),
.io_dataIn_1374(dataIn[1374]),
.io_dataIn_1375(dataIn[1375]),
.io_dataIn_1376(dataIn[1376]),
.io_dataIn_1377(dataIn[1377]),
.io_dataIn_1378(dataIn[1378]),
.io_dataIn_1379(dataIn[1379]),
.io_dataIn_1380(dataIn[1380]),
.io_dataIn_1381(dataIn[1381]),
.io_dataIn_1382(dataIn[1382]),
.io_dataIn_1383(dataIn[1383]),
.io_dataIn_1384(dataIn[1384]),
.io_dataIn_1385(dataIn[1385]),
.io_dataIn_1386(dataIn[1386]),
.io_dataIn_1387(dataIn[1387]),
.io_dataIn_1388(dataIn[1388]),
.io_dataIn_1389(dataIn[1389]),
.io_dataIn_1390(dataIn[1390]),
.io_dataIn_1391(dataIn[1391]),
.io_dataIn_1392(dataIn[1392]),
.io_dataIn_1393(dataIn[1393]),
.io_dataIn_1394(dataIn[1394]),
.io_dataIn_1395(dataIn[1395]),
.io_dataIn_1396(dataIn[1396]),
.io_dataIn_1397(dataIn[1397]),
.io_dataIn_1398(dataIn[1398]),
.io_dataIn_1399(dataIn[1399]),
.io_dataIn_1400(dataIn[1400]),
.io_dataIn_1401(dataIn[1401]),
.io_dataIn_1402(dataIn[1402]),
.io_dataIn_1403(dataIn[1403]),
.io_dataIn_1404(dataIn[1404]),
.io_dataIn_1405(dataIn[1405]),
.io_dataIn_1406(dataIn[1406]),
.io_dataIn_1407(dataIn[1407]),
.io_dataIn_1408(dataIn[1408]),
.io_dataIn_1409(dataIn[1409]),
.io_dataIn_1410(dataIn[1410]),
.io_dataIn_1411(dataIn[1411]),
.io_dataIn_1412(dataIn[1412]),
.io_dataIn_1413(dataIn[1413]),
.io_dataIn_1414(dataIn[1414]),
.io_dataIn_1415(dataIn[1415]),
.io_dataIn_1416(dataIn[1416]),
.io_dataIn_1417(dataIn[1417]),
.io_dataIn_1418(dataIn[1418]),
.io_dataIn_1419(dataIn[1419]),
.io_dataIn_1420(dataIn[1420]),
.io_dataIn_1421(dataIn[1421]),
.io_dataIn_1422(dataIn[1422]),
.io_dataIn_1423(dataIn[1423]),
.io_dataIn_1424(dataIn[1424]),
.io_dataIn_1425(dataIn[1425]),
.io_dataIn_1426(dataIn[1426]),
.io_dataIn_1427(dataIn[1427]),
.io_dataIn_1428(dataIn[1428]),
.io_dataIn_1429(dataIn[1429]),
.io_dataIn_1430(dataIn[1430]),
.io_dataIn_1431(dataIn[1431]),
.io_dataIn_1432(dataIn[1432]),
.io_dataIn_1433(dataIn[1433]),
.io_dataIn_1434(dataIn[1434]),
.io_dataIn_1435(dataIn[1435]),
.io_dataIn_1436(dataIn[1436]),
.io_dataIn_1437(dataIn[1437]),
.io_dataIn_1438(dataIn[1438]),
.io_dataIn_1439(dataIn[1439]),
.io_dataIn_1440(dataIn[1440]),
.io_dataIn_1441(dataIn[1441]),
.io_dataIn_1442(dataIn[1442]),
.io_dataIn_1443(dataIn[1443]),
.io_dataIn_1444(dataIn[1444]),
.io_dataIn_1445(dataIn[1445]),
.io_dataIn_1446(dataIn[1446]),
.io_dataIn_1447(dataIn[1447]),
.io_dataIn_1448(dataIn[1448]),
.io_dataIn_1449(dataIn[1449]),
.io_dataIn_1450(dataIn[1450]),
.io_dataIn_1451(dataIn[1451]),
.io_dataIn_1452(dataIn[1452]),
.io_dataIn_1453(dataIn[1453]),
.io_dataIn_1454(dataIn[1454]),
.io_dataIn_1455(dataIn[1455]),
.io_dataIn_1456(dataIn[1456]),
.io_dataIn_1457(dataIn[1457]),
.io_dataIn_1458(dataIn[1458]),
.io_dataIn_1459(dataIn[1459]),
.io_dataIn_1460(dataIn[1460]),
.io_dataIn_1461(dataIn[1461]),
.io_dataIn_1462(dataIn[1462]),
.io_dataIn_1463(dataIn[1463]),
.io_dataIn_1464(dataIn[1464]),
.io_dataIn_1465(dataIn[1465]),
.io_dataIn_1466(dataIn[1466]),
.io_dataIn_1467(dataIn[1467]),
.io_dataIn_1468(dataIn[1468]),
.io_dataIn_1469(dataIn[1469]),
.io_dataIn_1470(dataIn[1470]),
.io_dataIn_1471(dataIn[1471]),
.io_dataIn_1472(dataIn[1472]),
.io_dataIn_1473(dataIn[1473]),
.io_dataIn_1474(dataIn[1474]),
.io_dataIn_1475(dataIn[1475]),
.io_dataIn_1476(dataIn[1476]),
.io_dataIn_1477(dataIn[1477]),
.io_dataIn_1478(dataIn[1478]),
.io_dataIn_1479(dataIn[1479]),
.io_dataIn_1480(dataIn[1480]),
.io_dataIn_1481(dataIn[1481]),
.io_dataIn_1482(dataIn[1482]),
.io_dataIn_1483(dataIn[1483]),
.io_dataIn_1484(dataIn[1484]),
.io_dataIn_1485(dataIn[1485]),
.io_dataIn_1486(dataIn[1486]),
.io_dataIn_1487(dataIn[1487]),
.io_dataIn_1488(dataIn[1488]),
.io_dataIn_1489(dataIn[1489]),
.io_dataIn_1490(dataIn[1490]),
.io_dataIn_1491(dataIn[1491]),
.io_dataIn_1492(dataIn[1492]),
.io_dataIn_1493(dataIn[1493]),
.io_dataIn_1494(dataIn[1494]),
.io_dataIn_1495(dataIn[1495]),
.io_dataIn_1496(dataIn[1496]),
.io_dataIn_1497(dataIn[1497]),
.io_dataIn_1498(dataIn[1498]),
.io_dataIn_1499(dataIn[1499]),
.io_dataIn_1500(dataIn[1500]),
.io_dataIn_1501(dataIn[1501]),
.io_dataIn_1502(dataIn[1502]),
.io_dataIn_1503(dataIn[1503]),
.io_dataIn_1504(dataIn[1504]),
.io_dataIn_1505(dataIn[1505]),
.io_dataIn_1506(dataIn[1506]),
.io_dataIn_1507(dataIn[1507]),
.io_dataIn_1508(dataIn[1508]),
.io_dataIn_1509(dataIn[1509]),
.io_dataIn_1510(dataIn[1510]),
.io_dataIn_1511(dataIn[1511]),
.io_dataIn_1512(dataIn[1512]),
.io_dataIn_1513(dataIn[1513]),
.io_dataIn_1514(dataIn[1514]),
.io_dataIn_1515(dataIn[1515]),
.io_dataIn_1516(dataIn[1516]),
.io_dataIn_1517(dataIn[1517]),
.io_dataIn_1518(dataIn[1518]),
.io_dataIn_1519(dataIn[1519]),
.io_dataIn_1520(dataIn[1520]),
.io_dataIn_1521(dataIn[1521]),
.io_dataIn_1522(dataIn[1522]),
.io_dataIn_1523(dataIn[1523]),
.io_dataIn_1524(dataIn[1524]),
.io_dataIn_1525(dataIn[1525]),
.io_dataIn_1526(dataIn[1526]),
.io_dataIn_1527(dataIn[1527]),
.io_dataIn_1528(dataIn[1528]),
.io_dataIn_1529(dataIn[1529]),
.io_dataIn_1530(dataIn[1530]),
.io_dataIn_1531(dataIn[1531]),
.io_dataIn_1532(dataIn[1532]),
.io_dataIn_1533(dataIn[1533]),
.io_dataIn_1534(dataIn[1534]),
.io_dataIn_1535(dataIn[1535]),
.io_dataIn_1536(dataIn[1536]),
.io_dataIn_1537(dataIn[1537]),
.io_dataIn_1538(dataIn[1538]),
.io_dataIn_1539(dataIn[1539]),
.io_dataIn_1540(dataIn[1540]),
.io_dataIn_1541(dataIn[1541]),
.io_dataIn_1542(dataIn[1542]),
.io_dataIn_1543(dataIn[1543]),
.io_dataIn_1544(dataIn[1544]),
.io_dataIn_1545(dataIn[1545]),
.io_dataIn_1546(dataIn[1546]),
.io_dataIn_1547(dataIn[1547]),
.io_dataIn_1548(dataIn[1548]),
.io_dataIn_1549(dataIn[1549]),
.io_dataIn_1550(dataIn[1550]),
.io_dataIn_1551(dataIn[1551]),
.io_dataIn_1552(dataIn[1552]),
.io_dataIn_1553(dataIn[1553]),
.io_dataIn_1554(dataIn[1554]),
.io_dataIn_1555(dataIn[1555]),
.io_dataIn_1556(dataIn[1556]),
.io_dataIn_1557(dataIn[1557]),
.io_dataIn_1558(dataIn[1558]),
.io_dataIn_1559(dataIn[1559]),
.io_dataIn_1560(dataIn[1560]),
.io_dataIn_1561(dataIn[1561]),
.io_dataIn_1562(dataIn[1562]),
.io_dataIn_1563(dataIn[1563]),
.io_dataIn_1564(dataIn[1564]),
.io_dataIn_1565(dataIn[1565]),
.io_dataIn_1566(dataIn[1566]),
.io_dataIn_1567(dataIn[1567]),
.io_dataIn_1568(dataIn[1568]),
.io_dataIn_1569(dataIn[1569]),
.io_dataIn_1570(dataIn[1570]),
.io_dataIn_1571(dataIn[1571]),
.io_dataIn_1572(dataIn[1572]),
.io_dataIn_1573(dataIn[1573]),
.io_dataIn_1574(dataIn[1574]),
.io_dataIn_1575(dataIn[1575]),
.io_dataIn_1576(dataIn[1576]),
.io_dataIn_1577(dataIn[1577]),
.io_dataIn_1578(dataIn[1578]),
.io_dataIn_1579(dataIn[1579]),
.io_dataIn_1580(dataIn[1580]),
.io_dataIn_1581(dataIn[1581]),
.io_dataIn_1582(dataIn[1582]),
.io_dataIn_1583(dataIn[1583]),
.io_dataIn_1584(dataIn[1584]),
.io_dataIn_1585(dataIn[1585]),
.io_dataIn_1586(dataIn[1586]),
.io_dataIn_1587(dataIn[1587]),
.io_dataIn_1588(dataIn[1588]),
.io_dataIn_1589(dataIn[1589]),
.io_dataIn_1590(dataIn[1590]),
.io_dataIn_1591(dataIn[1591]),
.io_dataIn_1592(dataIn[1592]),
.io_dataIn_1593(dataIn[1593]),
.io_dataIn_1594(dataIn[1594]),
.io_dataIn_1595(dataIn[1595]),
.io_dataIn_1596(dataIn[1596]),
.io_dataIn_1597(dataIn[1597]),
.io_dataIn_1598(dataIn[1598]),
.io_dataIn_1599(dataIn[1599]),
.io_dataIn_1600(dataIn[1600]),
.io_dataIn_1601(dataIn[1601]),
.io_dataIn_1602(dataIn[1602]),
.io_dataIn_1603(dataIn[1603]),
.io_dataIn_1604(dataIn[1604]),
.io_dataIn_1605(dataIn[1605]),
.io_dataIn_1606(dataIn[1606]),
.io_dataIn_1607(dataIn[1607]),
.io_dataIn_1608(dataIn[1608]),
.io_dataIn_1609(dataIn[1609]),
.io_dataIn_1610(dataIn[1610]),
.io_dataIn_1611(dataIn[1611]),
.io_dataIn_1612(dataIn[1612]),
.io_dataIn_1613(dataIn[1613]),
.io_dataIn_1614(dataIn[1614]),
.io_dataIn_1615(dataIn[1615]),
.io_dataIn_1616(dataIn[1616]),
.io_dataIn_1617(dataIn[1617]),
.io_dataIn_1618(dataIn[1618]),
.io_dataIn_1619(dataIn[1619]),
.io_dataIn_1620(dataIn[1620]),
.io_dataIn_1621(dataIn[1621]),
.io_dataIn_1622(dataIn[1622]),
.io_dataIn_1623(dataIn[1623]),
.io_dataIn_1624(dataIn[1624]),
.io_dataIn_1625(dataIn[1625]),
.io_dataIn_1626(dataIn[1626]),
.io_dataIn_1627(dataIn[1627]),
.io_dataIn_1628(dataIn[1628]),
.io_dataIn_1629(dataIn[1629]),
.io_dataIn_1630(dataIn[1630]),
.io_dataIn_1631(dataIn[1631]),
.io_dataIn_1632(dataIn[1632]),
.io_dataIn_1633(dataIn[1633]),
.io_dataIn_1634(dataIn[1634]),
.io_dataIn_1635(dataIn[1635]),
.io_dataIn_1636(dataIn[1636]),
.io_dataIn_1637(dataIn[1637]),
.io_dataIn_1638(dataIn[1638]),
.io_dataIn_1639(dataIn[1639]),
.io_dataIn_1640(dataIn[1640]),
.io_dataIn_1641(dataIn[1641]),
.io_dataIn_1642(dataIn[1642]),
.io_dataIn_1643(dataIn[1643]),
.io_dataIn_1644(dataIn[1644]),
.io_dataIn_1645(dataIn[1645]),
.io_dataIn_1646(dataIn[1646]),
.io_dataIn_1647(dataIn[1647]),
.io_dataIn_1648(dataIn[1648]),
.io_dataIn_1649(dataIn[1649]),
.io_dataIn_1650(dataIn[1650]),
.io_dataIn_1651(dataIn[1651]),
.io_dataIn_1652(dataIn[1652]),
.io_dataIn_1653(dataIn[1653]),
.io_dataIn_1654(dataIn[1654]),
.io_dataIn_1655(dataIn[1655]),
.io_dataIn_1656(dataIn[1656]),
.io_dataIn_1657(dataIn[1657]),
.io_dataIn_1658(dataIn[1658]),
.io_dataIn_1659(dataIn[1659]),
.io_dataIn_1660(dataIn[1660]),
.io_dataIn_1661(dataIn[1661]),
.io_dataIn_1662(dataIn[1662]),
.io_dataIn_1663(dataIn[1663]),
.io_dataIn_1664(dataIn[1664]),
.io_dataIn_1665(dataIn[1665]),
.io_dataIn_1666(dataIn[1666]),
.io_dataIn_1667(dataIn[1667]),
.io_dataIn_1668(dataIn[1668]),
.io_dataIn_1669(dataIn[1669]),
.io_dataIn_1670(dataIn[1670]),
.io_dataIn_1671(dataIn[1671]),
.io_dataIn_1672(dataIn[1672]),
.io_dataIn_1673(dataIn[1673]),
.io_dataIn_1674(dataIn[1674]),
.io_dataIn_1675(dataIn[1675]),
.io_dataIn_1676(dataIn[1676]),
.io_dataIn_1677(dataIn[1677]),
.io_dataIn_1678(dataIn[1678]),
.io_dataIn_1679(dataIn[1679]),
.io_dataIn_1680(dataIn[1680]),
.io_dataIn_1681(dataIn[1681]),
.io_dataIn_1682(dataIn[1682]),
.io_dataIn_1683(dataIn[1683]),
.io_dataIn_1684(dataIn[1684]),
.io_dataIn_1685(dataIn[1685]),
.io_dataIn_1686(dataIn[1686]),
.io_dataIn_1687(dataIn[1687]),
.io_dataIn_1688(dataIn[1688]),
.io_dataIn_1689(dataIn[1689]),
.io_dataIn_1690(dataIn[1690]),
.io_dataIn_1691(dataIn[1691]),
.io_dataIn_1692(dataIn[1692]),
.io_dataIn_1693(dataIn[1693]),
.io_dataIn_1694(dataIn[1694]),
.io_dataIn_1695(dataIn[1695]),
.io_dataIn_1696(dataIn[1696]),
.io_dataIn_1697(dataIn[1697]),
.io_dataIn_1698(dataIn[1698]),
.io_dataIn_1699(dataIn[1699]),
.io_dataIn_1700(dataIn[1700]),
.io_dataIn_1701(dataIn[1701]),
.io_dataIn_1702(dataIn[1702]),
.io_dataIn_1703(dataIn[1703]),
.io_dataIn_1704(dataIn[1704]),
.io_dataIn_1705(dataIn[1705]),
.io_dataIn_1706(dataIn[1706]),
.io_dataIn_1707(dataIn[1707]),
.io_dataIn_1708(dataIn[1708]),
.io_dataIn_1709(dataIn[1709]),
.io_dataIn_1710(dataIn[1710]),
.io_dataIn_1711(dataIn[1711]),
.io_dataIn_1712(dataIn[1712]),
.io_dataIn_1713(dataIn[1713]),
.io_dataIn_1714(dataIn[1714]),
.io_dataIn_1715(dataIn[1715]),
.io_dataIn_1716(dataIn[1716]),
.io_dataIn_1717(dataIn[1717]),
.io_dataIn_1718(dataIn[1718]),
.io_dataIn_1719(dataIn[1719]),
.io_dataIn_1720(dataIn[1720]),
.io_dataIn_1721(dataIn[1721]),
.io_dataIn_1722(dataIn[1722]),
.io_dataIn_1723(dataIn[1723]),
.io_dataIn_1724(dataIn[1724]),
.io_dataIn_1725(dataIn[1725]),
.io_dataIn_1726(dataIn[1726]),
.io_dataIn_1727(dataIn[1727]),
.io_dataIn_1728(dataIn[1728]),
.io_dataIn_1729(dataIn[1729]),
.io_dataIn_1730(dataIn[1730]),
.io_dataIn_1731(dataIn[1731]),
.io_dataIn_1732(dataIn[1732]),
.io_dataIn_1733(dataIn[1733]),
.io_dataIn_1734(dataIn[1734]),
.io_dataIn_1735(dataIn[1735]),
.io_dataIn_1736(dataIn[1736]),
.io_dataIn_1737(dataIn[1737]),
.io_dataIn_1738(dataIn[1738]),
.io_dataIn_1739(dataIn[1739]),
.io_dataIn_1740(dataIn[1740]),
.io_dataIn_1741(dataIn[1741]),
.io_dataIn_1742(dataIn[1742]),
.io_dataIn_1743(dataIn[1743]),
.io_dataIn_1744(dataIn[1744]),
.io_dataIn_1745(dataIn[1745]),
.io_dataIn_1746(dataIn[1746]),
.io_dataIn_1747(dataIn[1747]),
.io_dataIn_1748(dataIn[1748]),
.io_dataIn_1749(dataIn[1749]),
.io_dataIn_1750(dataIn[1750]),
.io_dataIn_1751(dataIn[1751]),
.io_dataIn_1752(dataIn[1752]),
.io_dataIn_1753(dataIn[1753]),
.io_dataIn_1754(dataIn[1754]),
.io_dataIn_1755(dataIn[1755]),
.io_dataIn_1756(dataIn[1756]),
.io_dataIn_1757(dataIn[1757]),
.io_dataIn_1758(dataIn[1758]),
.io_dataIn_1759(dataIn[1759]),
.io_dataIn_1760(dataIn[1760]),
.io_dataIn_1761(dataIn[1761]),
.io_dataIn_1762(dataIn[1762]),
.io_dataIn_1763(dataIn[1763]),
.io_dataIn_1764(dataIn[1764]),
.io_dataIn_1765(dataIn[1765]),
.io_dataIn_1766(dataIn[1766]),
.io_dataIn_1767(dataIn[1767]),
.io_dataIn_1768(dataIn[1768]),
.io_dataIn_1769(dataIn[1769]),
.io_dataIn_1770(dataIn[1770]),
.io_dataIn_1771(dataIn[1771]),
.io_dataIn_1772(dataIn[1772]),
.io_dataIn_1773(dataIn[1773]),
.io_dataIn_1774(dataIn[1774]),
.io_dataIn_1775(dataIn[1775]),
.io_dataIn_1776(dataIn[1776]),
.io_dataIn_1777(dataIn[1777]),
.io_dataIn_1778(dataIn[1778]),
.io_dataIn_1779(dataIn[1779]),
.io_dataIn_1780(dataIn[1780]),
.io_dataIn_1781(dataIn[1781]),
.io_dataIn_1782(dataIn[1782]),
.io_dataIn_1783(dataIn[1783]),
.io_dataIn_1784(dataIn[1784]),
.io_dataIn_1785(dataIn[1785]),
.io_dataIn_1786(dataIn[1786]),
.io_dataIn_1787(dataIn[1787]),
.io_dataIn_1788(dataIn[1788]),
.io_dataIn_1789(dataIn[1789]),
.io_dataIn_1790(dataIn[1790]),
.io_dataIn_1791(dataIn[1791]),
.io_dataIn_1792(dataIn[1792]),
.io_dataIn_1793(dataIn[1793]),
.io_dataIn_1794(dataIn[1794]),
.io_dataIn_1795(dataIn[1795]),
.io_dataIn_1796(dataIn[1796]),
.io_dataIn_1797(dataIn[1797]),
.io_dataIn_1798(dataIn[1798]),
.io_dataIn_1799(dataIn[1799]),
.io_dataIn_1800(dataIn[1800]),
.io_dataIn_1801(dataIn[1801]),
.io_dataIn_1802(dataIn[1802]),
.io_dataIn_1803(dataIn[1803]),
.io_dataIn_1804(dataIn[1804]),
.io_dataIn_1805(dataIn[1805]),
.io_dataIn_1806(dataIn[1806]),
.io_dataIn_1807(dataIn[1807]),
.io_dataIn_1808(dataIn[1808]),
.io_dataIn_1809(dataIn[1809]),
.io_dataIn_1810(dataIn[1810]),
.io_dataIn_1811(dataIn[1811]),
.io_dataIn_1812(dataIn[1812]),
.io_dataIn_1813(dataIn[1813]),
.io_dataIn_1814(dataIn[1814]),
.io_dataIn_1815(dataIn[1815]),
.io_dataIn_1816(dataIn[1816]),
.io_dataIn_1817(dataIn[1817]),
.io_dataIn_1818(dataIn[1818]),
.io_dataIn_1819(dataIn[1819]),
.io_dataIn_1820(dataIn[1820]),
.io_dataIn_1821(dataIn[1821]),
.io_dataIn_1822(dataIn[1822]),
.io_dataIn_1823(dataIn[1823]),
.io_dataIn_1824(dataIn[1824]),
.io_dataIn_1825(dataIn[1825]),
.io_dataIn_1826(dataIn[1826]),
.io_dataIn_1827(dataIn[1827]),
.io_dataIn_1828(dataIn[1828]),
.io_dataIn_1829(dataIn[1829]),
.io_dataIn_1830(dataIn[1830]),
.io_dataIn_1831(dataIn[1831]),
.io_dataIn_1832(dataIn[1832]),
.io_dataIn_1833(dataIn[1833]),
.io_dataIn_1834(dataIn[1834]),
.io_dataIn_1835(dataIn[1835]),
.io_dataIn_1836(dataIn[1836]),
.io_dataIn_1837(dataIn[1837]),
.io_dataIn_1838(dataIn[1838]),
.io_dataIn_1839(dataIn[1839]),
.io_dataIn_1840(dataIn[1840]),
.io_dataIn_1841(dataIn[1841]),
.io_dataIn_1842(dataIn[1842]),
.io_dataIn_1843(dataIn[1843]),
.io_dataIn_1844(dataIn[1844]),
.io_dataIn_1845(dataIn[1845]),
.io_dataIn_1846(dataIn[1846]),
.io_dataIn_1847(dataIn[1847]),
.io_dataIn_1848(dataIn[1848]),
.io_dataIn_1849(dataIn[1849]),
.io_dataIn_1850(dataIn[1850]),
.io_dataIn_1851(dataIn[1851]),
.io_dataIn_1852(dataIn[1852]),
.io_dataIn_1853(dataIn[1853]),
.io_dataIn_1854(dataIn[1854]),
.io_dataIn_1855(dataIn[1855]),
.io_dataIn_1856(dataIn[1856]),
.io_dataIn_1857(dataIn[1857]),
.io_dataIn_1858(dataIn[1858]),
.io_dataIn_1859(dataIn[1859]),
.io_dataIn_1860(dataIn[1860]),
.io_dataIn_1861(dataIn[1861]),
.io_dataIn_1862(dataIn[1862]),
.io_dataIn_1863(dataIn[1863]),
.io_dataIn_1864(dataIn[1864]),
.io_dataIn_1865(dataIn[1865]),
.io_dataIn_1866(dataIn[1866]),
.io_dataIn_1867(dataIn[1867]),
.io_dataIn_1868(dataIn[1868]),
.io_dataIn_1869(dataIn[1869]),
.io_dataIn_1870(dataIn[1870]),
.io_dataIn_1871(dataIn[1871]),
.io_dataIn_1872(dataIn[1872]),
.io_dataIn_1873(dataIn[1873]),
.io_dataIn_1874(dataIn[1874]),
.io_dataIn_1875(dataIn[1875]),
.io_dataIn_1876(dataIn[1876]),
.io_dataIn_1877(dataIn[1877]),
.io_dataIn_1878(dataIn[1878]),
.io_dataIn_1879(dataIn[1879]),
.io_dataIn_1880(dataIn[1880]),
.io_dataIn_1881(dataIn[1881]),
.io_dataIn_1882(dataIn[1882]),
.io_dataIn_1883(dataIn[1883]),
.io_dataIn_1884(dataIn[1884]),
.io_dataIn_1885(dataIn[1885]),
.io_dataIn_1886(dataIn[1886]),
.io_dataIn_1887(dataIn[1887]),
.io_dataIn_1888(dataIn[1888]),
.io_dataIn_1889(dataIn[1889]),
.io_dataIn_1890(dataIn[1890]),
.io_dataIn_1891(dataIn[1891]),
.io_dataIn_1892(dataIn[1892]),
.io_dataIn_1893(dataIn[1893]),
.io_dataIn_1894(dataIn[1894]),
.io_dataIn_1895(dataIn[1895]),
.io_dataIn_1896(dataIn[1896]),
.io_dataIn_1897(dataIn[1897]),
.io_dataIn_1898(dataIn[1898]),
.io_dataIn_1899(dataIn[1899]),
.io_dataIn_1900(dataIn[1900]),
.io_dataIn_1901(dataIn[1901]),
.io_dataIn_1902(dataIn[1902]),
.io_dataIn_1903(dataIn[1903]),
.io_dataIn_1904(dataIn[1904]),
.io_dataIn_1905(dataIn[1905]),
.io_dataIn_1906(dataIn[1906]),
.io_dataIn_1907(dataIn[1907]),
.io_dataIn_1908(dataIn[1908]),
.io_dataIn_1909(dataIn[1909]),
.io_dataIn_1910(dataIn[1910]),
.io_dataIn_1911(dataIn[1911]),
.io_dataIn_1912(dataIn[1912]),
.io_dataIn_1913(dataIn[1913]),
.io_dataIn_1914(dataIn[1914]),
.io_dataIn_1915(dataIn[1915]),
.io_dataIn_1916(dataIn[1916]),
.io_dataIn_1917(dataIn[1917]),
.io_dataIn_1918(dataIn[1918]),
.io_dataIn_1919(dataIn[1919]),
.io_dataIn_1920(dataIn[1920]),
.io_dataIn_1921(dataIn[1921]),
.io_dataIn_1922(dataIn[1922]),
.io_dataIn_1923(dataIn[1923]),
.io_dataIn_1924(dataIn[1924]),
.io_dataIn_1925(dataIn[1925]),
.io_dataIn_1926(dataIn[1926]),
.io_dataIn_1927(dataIn[1927]),
.io_dataIn_1928(dataIn[1928]),
.io_dataIn_1929(dataIn[1929]),
.io_dataIn_1930(dataIn[1930]),
.io_dataIn_1931(dataIn[1931]),
.io_dataIn_1932(dataIn[1932]),
.io_dataIn_1933(dataIn[1933]),
.io_dataIn_1934(dataIn[1934]),
.io_dataIn_1935(dataIn[1935]),
.io_dataIn_1936(dataIn[1936]),
.io_dataIn_1937(dataIn[1937]),
.io_dataIn_1938(dataIn[1938]),
.io_dataIn_1939(dataIn[1939]),
.io_dataIn_1940(dataIn[1940]),
.io_dataIn_1941(dataIn[1941]),
.io_dataIn_1942(dataIn[1942]),
.io_dataIn_1943(dataIn[1943]),
.io_dataIn_1944(dataIn[1944]),
.io_dataIn_1945(dataIn[1945]),
.io_dataIn_1946(dataIn[1946]),
.io_dataIn_1947(dataIn[1947]),
.io_dataIn_1948(dataIn[1948]),
.io_dataIn_1949(dataIn[1949]),
.io_dataIn_1950(dataIn[1950]),
.io_dataIn_1951(dataIn[1951]),
.io_dataIn_1952(dataIn[1952]),
.io_dataIn_1953(dataIn[1953]),
.io_dataIn_1954(dataIn[1954]),
.io_dataIn_1955(dataIn[1955]),
.io_dataIn_1956(dataIn[1956]),
.io_dataIn_1957(dataIn[1957]),
.io_dataIn_1958(dataIn[1958]),
.io_dataIn_1959(dataIn[1959]),
.io_dataIn_1960(dataIn[1960]),
.io_dataIn_1961(dataIn[1961]),
.io_dataIn_1962(dataIn[1962]),
.io_dataIn_1963(dataIn[1963]),
.io_dataIn_1964(dataIn[1964]),
.io_dataIn_1965(dataIn[1965]),
.io_dataIn_1966(dataIn[1966]),
.io_dataIn_1967(dataIn[1967]),
.io_dataIn_1968(dataIn[1968]),
.io_dataIn_1969(dataIn[1969]),
.io_dataIn_1970(dataIn[1970]),
.io_dataIn_1971(dataIn[1971]),
.io_dataIn_1972(dataIn[1972]),
.io_dataIn_1973(dataIn[1973]),
.io_dataIn_1974(dataIn[1974]),
.io_dataIn_1975(dataIn[1975]),
.io_dataIn_1976(dataIn[1976]),
.io_dataIn_1977(dataIn[1977]),
.io_dataIn_1978(dataIn[1978]),
.io_dataIn_1979(dataIn[1979]),
.io_dataIn_1980(dataIn[1980]),
.io_dataIn_1981(dataIn[1981]),
.io_dataIn_1982(dataIn[1982]),
.io_dataIn_1983(dataIn[1983]),
.io_dataIn_1984(dataIn[1984]),
.io_dataIn_1985(dataIn[1985]),
.io_dataIn_1986(dataIn[1986]),
.io_dataIn_1987(dataIn[1987]),
.io_dataIn_1988(dataIn[1988]),
.io_dataIn_1989(dataIn[1989]),
.io_dataIn_1990(dataIn[1990]),
.io_dataIn_1991(dataIn[1991]),
.io_dataIn_1992(dataIn[1992]),
.io_dataIn_1993(dataIn[1993]),
.io_dataIn_1994(dataIn[1994]),
.io_dataIn_1995(dataIn[1995]),
.io_dataIn_1996(dataIn[1996]),
.io_dataIn_1997(dataIn[1997]),
.io_dataIn_1998(dataIn[1998]),
.io_dataIn_1999(dataIn[1999]),
.io_dataIn_2000(dataIn[2000]),
.io_dataIn_2001(dataIn[2001]),
.io_dataIn_2002(dataIn[2002]),
.io_dataIn_2003(dataIn[2003]),
.io_dataIn_2004(dataIn[2004]),
.io_dataIn_2005(dataIn[2005]),
.io_dataIn_2006(dataIn[2006]),
.io_dataIn_2007(dataIn[2007]),
.io_dataIn_2008(dataIn[2008]),
.io_dataIn_2009(dataIn[2009]),
.io_dataIn_2010(dataIn[2010]),
.io_dataIn_2011(dataIn[2011]),
.io_dataIn_2012(dataIn[2012]),
.io_dataIn_2013(dataIn[2013]),
.io_dataIn_2014(dataIn[2014]),
.io_dataIn_2015(dataIn[2015]),
.io_dataIn_2016(dataIn[2016]),
.io_dataIn_2017(dataIn[2017]),
.io_dataIn_2018(dataIn[2018]),
.io_dataIn_2019(dataIn[2019]),
.io_dataIn_2020(dataIn[2020]),
.io_dataIn_2021(dataIn[2021]),
.io_dataIn_2022(dataIn[2022]),
.io_dataIn_2023(dataIn[2023]),
.io_dataIn_2024(dataIn[2024]),
.io_dataIn_2025(dataIn[2025]),
.io_dataIn_2026(dataIn[2026]),
.io_dataIn_2027(dataIn[2027]),
.io_dataIn_2028(dataIn[2028]),
.io_dataIn_2029(dataIn[2029]),
.io_dataIn_2030(dataIn[2030]),
.io_dataIn_2031(dataIn[2031]),
.io_dataIn_2032(dataIn[2032]),
.io_dataIn_2033(dataIn[2033]),
.io_dataIn_2034(dataIn[2034]),
.io_dataIn_2035(dataIn[2035]),
.io_dataIn_2036(dataIn[2036]),
.io_dataIn_2037(dataIn[2037]),
.io_dataIn_2038(dataIn[2038]),
.io_dataIn_2039(dataIn[2039]),
.io_dataIn_2040(dataIn[2040]),
.io_dataIn_2041(dataIn[2041]),
.io_dataIn_2042(dataIn[2042]),
.io_dataIn_2043(dataIn[2043]),
.io_dataIn_2044(dataIn[2044]),
.io_dataIn_2045(dataIn[2045]),
.io_dataIn_2046(dataIn[2046]),
.io_dataIn_2047(dataIn[2047]),
.io_dataIn_2048(dataIn[2048]),
.io_dataIn_2049(dataIn[2049]),
.io_dataIn_2050(dataIn[2050]),
.io_dataIn_2051(dataIn[2051]),
.io_dataIn_2052(dataIn[2052]),
.io_dataIn_2053(dataIn[2053]),
.io_dataIn_2054(dataIn[2054]),
.io_dataIn_2055(dataIn[2055]),
.io_dataIn_2056(dataIn[2056]),
.io_dataIn_2057(dataIn[2057]),
.io_dataIn_2058(dataIn[2058]),
.io_dataIn_2059(dataIn[2059]),
.io_dataIn_2060(dataIn[2060]),
.io_dataIn_2061(dataIn[2061]),
.io_dataIn_2062(dataIn[2062]),
.io_dataIn_2063(dataIn[2063]),
.io_dataIn_2064(dataIn[2064]),
.io_dataIn_2065(dataIn[2065]),
.io_dataIn_2066(dataIn[2066]),
.io_dataIn_2067(dataIn[2067]),
.io_dataIn_2068(dataIn[2068]),
.io_dataIn_2069(dataIn[2069]),
.io_dataIn_2070(dataIn[2070]),
.io_dataIn_2071(dataIn[2071]),
.io_dataIn_2072(dataIn[2072]),
.io_dataIn_2073(dataIn[2073]),
.io_dataIn_2074(dataIn[2074]),
.io_dataIn_2075(dataIn[2075]),
.io_dataIn_2076(dataIn[2076]),
.io_dataIn_2077(dataIn[2077]),
.io_dataIn_2078(dataIn[2078]),
.io_dataIn_2079(dataIn[2079]),
.io_dataIn_2080(dataIn[2080]),
.io_dataIn_2081(dataIn[2081]),
.io_dataIn_2082(dataIn[2082]),
.io_dataIn_2083(dataIn[2083]),
.io_dataIn_2084(dataIn[2084]),
.io_dataIn_2085(dataIn[2085]),
.io_dataIn_2086(dataIn[2086]),
.io_dataIn_2087(dataIn[2087]),
.io_dataIn_2088(dataIn[2088]),
.io_dataIn_2089(dataIn[2089]),
.io_dataIn_2090(dataIn[2090]),
.io_dataIn_2091(dataIn[2091]),
.io_dataIn_2092(dataIn[2092]),
.io_dataIn_2093(dataIn[2093]),
.io_dataIn_2094(dataIn[2094]),
.io_dataIn_2095(dataIn[2095]),
.io_dataIn_2096(dataIn[2096]),
.io_dataIn_2097(dataIn[2097]),
.io_dataIn_2098(dataIn[2098]),
.io_dataIn_2099(dataIn[2099]),
.io_dataIn_2100(dataIn[2100]),
.io_dataIn_2101(dataIn[2101]),
.io_dataIn_2102(dataIn[2102]),
.io_dataIn_2103(dataIn[2103]),
.io_dataIn_2104(dataIn[2104]),
.io_dataIn_2105(dataIn[2105]),
.io_dataIn_2106(dataIn[2106]),
.io_dataIn_2107(dataIn[2107]),
.io_dataIn_2108(dataIn[2108]),
.io_dataIn_2109(dataIn[2109]),
.io_dataIn_2110(dataIn[2110]),
.io_dataIn_2111(dataIn[2111]),
.io_dataIn_2112(dataIn[2112]),
.io_dataIn_2113(dataIn[2113]),
.io_dataIn_2114(dataIn[2114]),
.io_dataIn_2115(dataIn[2115]),
.io_dataIn_2116(dataIn[2116]),
.io_dataIn_2117(dataIn[2117]),
.io_dataIn_2118(dataIn[2118]),
.io_dataIn_2119(dataIn[2119]),
.io_dataIn_2120(dataIn[2120]),
.io_dataIn_2121(dataIn[2121]),
.io_dataIn_2122(dataIn[2122]),
.io_dataIn_2123(dataIn[2123]),
.io_dataIn_2124(dataIn[2124]),
.io_dataIn_2125(dataIn[2125]),
.io_dataIn_2126(dataIn[2126]),
.io_dataIn_2127(dataIn[2127]),
.io_dataIn_2128(dataIn[2128]),
.io_dataIn_2129(dataIn[2129]),
.io_dataIn_2130(dataIn[2130]),
.io_dataIn_2131(dataIn[2131]),
.io_dataIn_2132(dataIn[2132]),
.io_dataIn_2133(dataIn[2133]),
.io_dataIn_2134(dataIn[2134]),
.io_dataIn_2135(dataIn[2135]),
.io_dataIn_2136(dataIn[2136]),
.io_dataIn_2137(dataIn[2137]),
.io_dataIn_2138(dataIn[2138]),
.io_dataIn_2139(dataIn[2139]),
.io_dataIn_2140(dataIn[2140]),
.io_dataIn_2141(dataIn[2141]),
.io_dataIn_2142(dataIn[2142]),
.io_dataIn_2143(dataIn[2143]),
.io_dataIn_2144(dataIn[2144]),
.io_dataIn_2145(dataIn[2145]),
.io_dataIn_2146(dataIn[2146]),
.io_dataIn_2147(dataIn[2147]),
.io_dataIn_2148(dataIn[2148]),
.io_dataIn_2149(dataIn[2149]),
.io_dataIn_2150(dataIn[2150]),
.io_dataIn_2151(dataIn[2151]),
.io_dataIn_2152(dataIn[2152]),
.io_dataIn_2153(dataIn[2153]),
.io_dataIn_2154(dataIn[2154]),
.io_dataIn_2155(dataIn[2155]),
.io_dataIn_2156(dataIn[2156]),
.io_dataIn_2157(dataIn[2157]),
.io_dataIn_2158(dataIn[2158]),
.io_dataIn_2159(dataIn[2159]),
.io_dataIn_2160(dataIn[2160]),
.io_dataIn_2161(dataIn[2161]),
.io_dataIn_2162(dataIn[2162]),
.io_dataIn_2163(dataIn[2163]),
.io_dataIn_2164(dataIn[2164]),
.io_dataIn_2165(dataIn[2165]),
.io_dataIn_2166(dataIn[2166]),
.io_dataIn_2167(dataIn[2167]),
.io_dataIn_2168(dataIn[2168]),
.io_dataIn_2169(dataIn[2169]),
.io_dataIn_2170(dataIn[2170]),
.io_dataIn_2171(dataIn[2171]),
.io_dataIn_2172(dataIn[2172]),
.io_dataIn_2173(dataIn[2173]),
.io_dataIn_2174(dataIn[2174]),
.io_dataIn_2175(dataIn[2175]),
.io_dataIn_2176(dataIn[2176]),
.io_dataIn_2177(dataIn[2177]),
.io_dataIn_2178(dataIn[2178]),
.io_dataIn_2179(dataIn[2179]),
.io_dataIn_2180(dataIn[2180]),
.io_dataIn_2181(dataIn[2181]),
.io_dataIn_2182(dataIn[2182]),
.io_dataIn_2183(dataIn[2183]),
.io_dataIn_2184(dataIn[2184]),
.io_dataIn_2185(dataIn[2185]),
.io_dataIn_2186(dataIn[2186]),
.io_dataIn_2187(dataIn[2187]),
.io_dataIn_2188(dataIn[2188]),
.io_dataIn_2189(dataIn[2189]),
.io_dataIn_2190(dataIn[2190]),
.io_dataIn_2191(dataIn[2191]),
.io_dataIn_2192(dataIn[2192]),
.io_dataIn_2193(dataIn[2193]),
.io_dataIn_2194(dataIn[2194]),
.io_dataIn_2195(dataIn[2195]),
.io_dataIn_2196(dataIn[2196]),
.io_dataIn_2197(dataIn[2197]),
.io_dataIn_2198(dataIn[2198]),
.io_dataIn_2199(dataIn[2199]),
.io_dataIn_2200(dataIn[2200]),
.io_dataIn_2201(dataIn[2201]),
.io_dataIn_2202(dataIn[2202]),
.io_dataIn_2203(dataIn[2203]),
.io_dataIn_2204(dataIn[2204]),
.io_dataIn_2205(dataIn[2205]),
.io_dataIn_2206(dataIn[2206]),
.io_dataIn_2207(dataIn[2207]),
.io_dataIn_2208(dataIn[2208]),
.io_dataIn_2209(dataIn[2209]),
.io_dataIn_2210(dataIn[2210]),
.io_dataIn_2211(dataIn[2211]),
.io_dataIn_2212(dataIn[2212]),
.io_dataIn_2213(dataIn[2213]),
.io_dataIn_2214(dataIn[2214]),
.io_dataIn_2215(dataIn[2215]),
.io_dataIn_2216(dataIn[2216]),
.io_dataIn_2217(dataIn[2217]),
.io_dataIn_2218(dataIn[2218]),
.io_dataIn_2219(dataIn[2219]),
.io_dataIn_2220(dataIn[2220]),
.io_dataIn_2221(dataIn[2221]),
.io_dataIn_2222(dataIn[2222]),
.io_dataIn_2223(dataIn[2223]),
.io_dataIn_2224(dataIn[2224]),
.io_dataIn_2225(dataIn[2225]),
.io_dataIn_2226(dataIn[2226]),
.io_dataIn_2227(dataIn[2227]),
.io_dataIn_2228(dataIn[2228]),
.io_dataIn_2229(dataIn[2229]),
.io_dataIn_2230(dataIn[2230]),
.io_dataIn_2231(dataIn[2231]),
.io_dataIn_2232(dataIn[2232]),
.io_dataIn_2233(dataIn[2233]),
.io_dataIn_2234(dataIn[2234]),
.io_dataIn_2235(dataIn[2235]),
.io_dataIn_2236(dataIn[2236]),
.io_dataIn_2237(dataIn[2237]),
.io_dataIn_2238(dataIn[2238]),
.io_dataIn_2239(dataIn[2239]),
.io_dataIn_2240(dataIn[2240]),
.io_dataIn_2241(dataIn[2241]),
.io_dataIn_2242(dataIn[2242]),
.io_dataIn_2243(dataIn[2243]),
.io_dataIn_2244(dataIn[2244]),
.io_dataIn_2245(dataIn[2245]),
.io_dataIn_2246(dataIn[2246]),
.io_dataIn_2247(dataIn[2247]),
.io_dataIn_2248(dataIn[2248]),
.io_dataIn_2249(dataIn[2249]),
.io_dataIn_2250(dataIn[2250]),
.io_dataIn_2251(dataIn[2251]),
.io_dataIn_2252(dataIn[2252]),
.io_dataIn_2253(dataIn[2253]),
.io_dataIn_2254(dataIn[2254]),
.io_dataIn_2255(dataIn[2255]),
.io_dataIn_2256(dataIn[2256]),
.io_dataIn_2257(dataIn[2257]),
.io_dataIn_2258(dataIn[2258]),
.io_dataIn_2259(dataIn[2259]),
.io_dataIn_2260(dataIn[2260]),
.io_dataIn_2261(dataIn[2261]),
.io_dataIn_2262(dataIn[2262]),
.io_dataIn_2263(dataIn[2263]),
.io_dataIn_2264(dataIn[2264]),
.io_dataIn_2265(dataIn[2265]),
.io_dataIn_2266(dataIn[2266]),
.io_dataIn_2267(dataIn[2267]),
.io_dataIn_2268(dataIn[2268]),
.io_dataIn_2269(dataIn[2269]),
.io_dataIn_2270(dataIn[2270]),
.io_dataIn_2271(dataIn[2271]),
.io_dataIn_2272(dataIn[2272]),
.io_dataIn_2273(dataIn[2273]),
.io_dataIn_2274(dataIn[2274]),
.io_dataIn_2275(dataIn[2275]),
.io_dataIn_2276(dataIn[2276]),
.io_dataIn_2277(dataIn[2277]),
.io_dataIn_2278(dataIn[2278]),
.io_dataIn_2279(dataIn[2279]),
.io_dataIn_2280(dataIn[2280]),
.io_dataIn_2281(dataIn[2281]),
.io_dataIn_2282(dataIn[2282]),
.io_dataIn_2283(dataIn[2283]),
.io_dataIn_2284(dataIn[2284]),
.io_dataIn_2285(dataIn[2285]),
.io_dataIn_2286(dataIn[2286]),
.io_dataIn_2287(dataIn[2287]),
.io_dataIn_2288(dataIn[2288]),
.io_dataIn_2289(dataIn[2289]),
.io_dataIn_2290(dataIn[2290]),
.io_dataIn_2291(dataIn[2291]),
.io_dataIn_2292(dataIn[2292]),
.io_dataIn_2293(dataIn[2293]),
.io_dataIn_2294(dataIn[2294]),
.io_dataIn_2295(dataIn[2295]),
.io_dataIn_2296(dataIn[2296]),
.io_dataIn_2297(dataIn[2297]),
.io_dataIn_2298(dataIn[2298]),
.io_dataIn_2299(dataIn[2299]),
.io_dataIn_2300(dataIn[2300]),
.io_dataIn_2301(dataIn[2301]),
.io_dataIn_2302(dataIn[2302]),
.io_dataIn_2303(dataIn[2303]),
.io_dataIn_2304(dataIn[2304]),
.io_dataIn_2305(dataIn[2305]),
.io_dataIn_2306(dataIn[2306]),
.io_dataIn_2307(dataIn[2307]),
.io_dataIn_2308(dataIn[2308]),
.io_dataIn_2309(dataIn[2309]),
.io_dataIn_2310(dataIn[2310]),
.io_dataIn_2311(dataIn[2311]),
.io_dataIn_2312(dataIn[2312]),
.io_dataIn_2313(dataIn[2313]),
.io_dataIn_2314(dataIn[2314]),
.io_dataIn_2315(dataIn[2315]),
.io_dataIn_2316(dataIn[2316]),
.io_dataIn_2317(dataIn[2317]),
.io_dataIn_2318(dataIn[2318]),
.io_dataIn_2319(dataIn[2319]),
.io_dataIn_2320(dataIn[2320]),
.io_dataIn_2321(dataIn[2321]),
.io_dataIn_2322(dataIn[2322]),
.io_dataIn_2323(dataIn[2323]),
.io_dataIn_2324(dataIn[2324]),
.io_dataIn_2325(dataIn[2325]),
.io_dataIn_2326(dataIn[2326]),
.io_dataIn_2327(dataIn[2327]),
.io_dataIn_2328(dataIn[2328]),
.io_dataIn_2329(dataIn[2329]),
.io_dataIn_2330(dataIn[2330]),
.io_dataIn_2331(dataIn[2331]),
.io_dataIn_2332(dataIn[2332]),
.io_dataIn_2333(dataIn[2333]),
.io_dataIn_2334(dataIn[2334]),
.io_dataIn_2335(dataIn[2335]),
.io_dataIn_2336(dataIn[2336]),
.io_dataIn_2337(dataIn[2337]),
.io_dataIn_2338(dataIn[2338]),
.io_dataIn_2339(dataIn[2339]),
.io_dataIn_2340(dataIn[2340]),
.io_dataIn_2341(dataIn[2341]),
.io_dataIn_2342(dataIn[2342]),
.io_dataIn_2343(dataIn[2343]),
.io_dataIn_2344(dataIn[2344]),
.io_dataIn_2345(dataIn[2345]),
.io_dataIn_2346(dataIn[2346]),
.io_dataIn_2347(dataIn[2347]),
.io_dataIn_2348(dataIn[2348]),
.io_dataIn_2349(dataIn[2349]),
.io_dataIn_2350(dataIn[2350]),
.io_dataIn_2351(dataIn[2351]),
.io_dataIn_2352(dataIn[2352]),
.io_dataIn_2353(dataIn[2353]),
.io_dataIn_2354(dataIn[2354]),
.io_dataIn_2355(dataIn[2355]),
.io_dataIn_2356(dataIn[2356]),
.io_dataIn_2357(dataIn[2357]),
.io_dataIn_2358(dataIn[2358]),
.io_dataIn_2359(dataIn[2359]),
.io_dataIn_2360(dataIn[2360]),
.io_dataIn_2361(dataIn[2361]),
.io_dataIn_2362(dataIn[2362]),
.io_dataIn_2363(dataIn[2363]),
.io_dataIn_2364(dataIn[2364]),
.io_dataIn_2365(dataIn[2365]),
.io_dataIn_2366(dataIn[2366]),
.io_dataIn_2367(dataIn[2367]),
.io_dataIn_2368(dataIn[2368]),
.io_dataIn_2369(dataIn[2369]),
.io_dataIn_2370(dataIn[2370]),
.io_dataIn_2371(dataIn[2371]),
.io_dataIn_2372(dataIn[2372]),
.io_dataIn_2373(dataIn[2373]),
.io_dataIn_2374(dataIn[2374]),
.io_dataIn_2375(dataIn[2375]),
.io_dataIn_2376(dataIn[2376]),
.io_dataIn_2377(dataIn[2377]),
.io_dataIn_2378(dataIn[2378]),
.io_dataIn_2379(dataIn[2379]),
.io_dataIn_2380(dataIn[2380]),
.io_dataIn_2381(dataIn[2381]),
.io_dataIn_2382(dataIn[2382]),
.io_dataIn_2383(dataIn[2383]),
.io_dataIn_2384(dataIn[2384]),
.io_dataIn_2385(dataIn[2385]),
.io_dataIn_2386(dataIn[2386]),
.io_dataIn_2387(dataIn[2387]),
.io_dataIn_2388(dataIn[2388]),
.io_dataIn_2389(dataIn[2389]),
.io_dataIn_2390(dataIn[2390]),
.io_dataIn_2391(dataIn[2391]),
.io_dataIn_2392(dataIn[2392]),
.io_dataIn_2393(dataIn[2393]),
.io_dataIn_2394(dataIn[2394]),
.io_dataIn_2395(dataIn[2395]),
.io_dataIn_2396(dataIn[2396]),
.io_dataIn_2397(dataIn[2397]),
.io_dataIn_2398(dataIn[2398]),
.io_dataIn_2399(dataIn[2399]),
.io_dataIn_2400(dataIn[2400]),
.io_dataIn_2401(dataIn[2401]),
.io_dataIn_2402(dataIn[2402]),
.io_dataIn_2403(dataIn[2403]),
.io_dataIn_2404(dataIn[2404]),
.io_dataIn_2405(dataIn[2405]),
.io_dataIn_2406(dataIn[2406]),
.io_dataIn_2407(dataIn[2407]),
.io_dataIn_2408(dataIn[2408]),
.io_dataIn_2409(dataIn[2409]),
.io_dataIn_2410(dataIn[2410]),
.io_dataIn_2411(dataIn[2411]),
.io_dataIn_2412(dataIn[2412]),
.io_dataIn_2413(dataIn[2413]),
.io_dataIn_2414(dataIn[2414]),
.io_dataIn_2415(dataIn[2415]),
.io_dataIn_2416(dataIn[2416]),
.io_dataIn_2417(dataIn[2417]),
.io_dataIn_2418(dataIn[2418]),
.io_dataIn_2419(dataIn[2419]),
.io_dataIn_2420(dataIn[2420]),
.io_dataIn_2421(dataIn[2421]),
.io_dataIn_2422(dataIn[2422]),
.io_dataIn_2423(dataIn[2423]),
.io_dataIn_2424(dataIn[2424]),
.io_dataIn_2425(dataIn[2425]),
.io_dataIn_2426(dataIn[2426]),
.io_dataIn_2427(dataIn[2427]),
.io_dataIn_2428(dataIn[2428]),
.io_dataIn_2429(dataIn[2429]),
.io_dataIn_2430(dataIn[2430]),
.io_dataIn_2431(dataIn[2431]),
.io_dataIn_2432(dataIn[2432]),
.io_dataIn_2433(dataIn[2433]),
.io_dataIn_2434(dataIn[2434]),
.io_dataIn_2435(dataIn[2435]),
.io_dataIn_2436(dataIn[2436]),
.io_dataIn_2437(dataIn[2437]),
.io_dataIn_2438(dataIn[2438]),
.io_dataIn_2439(dataIn[2439]),
.io_dataIn_2440(dataIn[2440]),
.io_dataIn_2441(dataIn[2441]),
.io_dataIn_2442(dataIn[2442]),
.io_dataIn_2443(dataIn[2443]),
.io_dataIn_2444(dataIn[2444]),
.io_dataIn_2445(dataIn[2445]),
.io_dataIn_2446(dataIn[2446]),
.io_dataIn_2447(dataIn[2447]),
.io_dataIn_2448(dataIn[2448]),
.io_dataIn_2449(dataIn[2449]),
.io_dataIn_2450(dataIn[2450]),
.io_dataIn_2451(dataIn[2451]),
.io_dataIn_2452(dataIn[2452]),
.io_dataIn_2453(dataIn[2453]),
.io_dataIn_2454(dataIn[2454]),
.io_dataIn_2455(dataIn[2455]),
.io_dataIn_2456(dataIn[2456]),
.io_dataIn_2457(dataIn[2457]),
.io_dataIn_2458(dataIn[2458]),
.io_dataIn_2459(dataIn[2459]),
.io_dataIn_2460(dataIn[2460]),
.io_dataIn_2461(dataIn[2461]),
.io_dataIn_2462(dataIn[2462]),
.io_dataIn_2463(dataIn[2463]),
.io_dataIn_2464(dataIn[2464]),
.io_dataIn_2465(dataIn[2465]),
.io_dataIn_2466(dataIn[2466]),
.io_dataIn_2467(dataIn[2467]),
.io_dataIn_2468(dataIn[2468]),
.io_dataIn_2469(dataIn[2469]),
.io_dataIn_2470(dataIn[2470]),
.io_dataIn_2471(dataIn[2471]),
.io_dataIn_2472(dataIn[2472]),
.io_dataIn_2473(dataIn[2473]),
.io_dataIn_2474(dataIn[2474]),
.io_dataIn_2475(dataIn[2475]),
.io_dataIn_2476(dataIn[2476]),
.io_dataIn_2477(dataIn[2477]),
.io_dataIn_2478(dataIn[2478]),
.io_dataIn_2479(dataIn[2479]),
.io_dataIn_2480(dataIn[2480]),
.io_dataIn_2481(dataIn[2481]),
.io_dataIn_2482(dataIn[2482]),
.io_dataIn_2483(dataIn[2483]),
.io_dataIn_2484(dataIn[2484]),
.io_dataIn_2485(dataIn[2485]),
.io_dataIn_2486(dataIn[2486]),
.io_dataIn_2487(dataIn[2487]),
.io_dataIn_2488(dataIn[2488]),
.io_dataIn_2489(dataIn[2489]),
.io_dataIn_2490(dataIn[2490]),
.io_dataIn_2491(dataIn[2491]),
.io_dataIn_2492(dataIn[2492]),
.io_dataIn_2493(dataIn[2493]),
.io_dataIn_2494(dataIn[2494]),
.io_dataIn_2495(dataIn[2495]),
.io_dataIn_2496(dataIn[2496]),
.io_dataIn_2497(dataIn[2497]),
.io_dataIn_2498(dataIn[2498]),
.io_dataIn_2499(dataIn[2499]),
.io_dataIn_2500(dataIn[2500]),
.io_dataIn_2501(dataIn[2501]),
.io_dataIn_2502(dataIn[2502]),
.io_dataIn_2503(dataIn[2503]),
.io_dataIn_2504(dataIn[2504]),
.io_dataIn_2505(dataIn[2505]),
.io_dataIn_2506(dataIn[2506]),
.io_dataIn_2507(dataIn[2507]),
.io_dataIn_2508(dataIn[2508]),
.io_dataIn_2509(dataIn[2509]),
.io_dataIn_2510(dataIn[2510]),
.io_dataIn_2511(dataIn[2511]),
.io_dataIn_2512(dataIn[2512]),
.io_dataIn_2513(dataIn[2513]),
.io_dataIn_2514(dataIn[2514]),
.io_dataIn_2515(dataIn[2515]),
.io_dataIn_2516(dataIn[2516]),
.io_dataIn_2517(dataIn[2517]),
.io_dataIn_2518(dataIn[2518]),
.io_dataIn_2519(dataIn[2519]),
.io_dataIn_2520(dataIn[2520]),
.io_dataIn_2521(dataIn[2521]),
.io_dataIn_2522(dataIn[2522]),
.io_dataIn_2523(dataIn[2523]),
.io_dataIn_2524(dataIn[2524]),
.io_dataIn_2525(dataIn[2525]),
.io_dataIn_2526(dataIn[2526]),
.io_dataIn_2527(dataIn[2527]),
.io_dataIn_2528(dataIn[2528]),
.io_dataIn_2529(dataIn[2529]),
.io_dataIn_2530(dataIn[2530]),
.io_dataIn_2531(dataIn[2531]),
.io_dataIn_2532(dataIn[2532]),
.io_dataIn_2533(dataIn[2533]),
.io_dataIn_2534(dataIn[2534]),
.io_dataIn_2535(dataIn[2535]),
.io_dataIn_2536(dataIn[2536]),
.io_dataIn_2537(dataIn[2537]),
.io_dataIn_2538(dataIn[2538]),
.io_dataIn_2539(dataIn[2539]),
.io_dataIn_2540(dataIn[2540]),
.io_dataIn_2541(dataIn[2541]),
.io_dataIn_2542(dataIn[2542]),
.io_dataIn_2543(dataIn[2543]),
.io_dataIn_2544(dataIn[2544]),
.io_dataIn_2545(dataIn[2545]),
.io_dataIn_2546(dataIn[2546]),
.io_dataIn_2547(dataIn[2547]),
.io_dataIn_2548(dataIn[2548]),
.io_dataIn_2549(dataIn[2549]),
.io_dataIn_2550(dataIn[2550]),
.io_dataIn_2551(dataIn[2551]),
.io_dataIn_2552(dataIn[2552]),
.io_dataIn_2553(dataIn[2553]),
.io_dataIn_2554(dataIn[2554]),
.io_dataIn_2555(dataIn[2555]),
.io_dataIn_2556(dataIn[2556]),
.io_dataIn_2557(dataIn[2557]),
.io_dataIn_2558(dataIn[2558]),
.io_dataIn_2559(dataIn[2559]),
.io_dataIn_2560(dataIn[2560]),
.io_dataIn_2561(dataIn[2561]),
.io_dataIn_2562(dataIn[2562]),
.io_dataIn_2563(dataIn[2563]),
.io_dataIn_2564(dataIn[2564]),
.io_dataIn_2565(dataIn[2565]),
.io_dataIn_2566(dataIn[2566]),
.io_dataIn_2567(dataIn[2567]),
.io_dataIn_2568(dataIn[2568]),
.io_dataIn_2569(dataIn[2569]),
.io_dataIn_2570(dataIn[2570]),
.io_dataIn_2571(dataIn[2571]),
.io_dataIn_2572(dataIn[2572]),
.io_dataIn_2573(dataIn[2573]),
.io_dataIn_2574(dataIn[2574]),
.io_dataIn_2575(dataIn[2575]),
.io_dataIn_2576(dataIn[2576]),
.io_dataIn_2577(dataIn[2577]),
.io_dataIn_2578(dataIn[2578]),
.io_dataIn_2579(dataIn[2579]),
.io_dataIn_2580(dataIn[2580]),
.io_dataIn_2581(dataIn[2581]),
.io_dataIn_2582(dataIn[2582]),
.io_dataIn_2583(dataIn[2583]),
.io_dataIn_2584(dataIn[2584]),
.io_dataIn_2585(dataIn[2585]),
.io_dataIn_2586(dataIn[2586]),
.io_dataIn_2587(dataIn[2587]),
.io_dataIn_2588(dataIn[2588]),
.io_dataIn_2589(dataIn[2589]),
.io_dataIn_2590(dataIn[2590]),
.io_dataIn_2591(dataIn[2591]),
.io_dataIn_2592(dataIn[2592]),
.io_dataIn_2593(dataIn[2593]),
.io_dataIn_2594(dataIn[2594]),
.io_dataIn_2595(dataIn[2595]),
.io_dataIn_2596(dataIn[2596]),
.io_dataIn_2597(dataIn[2597]),
.io_dataIn_2598(dataIn[2598]),
.io_dataIn_2599(dataIn[2599]),
.io_dataIn_2600(dataIn[2600]),
.io_dataIn_2601(dataIn[2601]),
.io_dataIn_2602(dataIn[2602]),
.io_dataIn_2603(dataIn[2603]),
.io_dataIn_2604(dataIn[2604]),
.io_dataIn_2605(dataIn[2605]),
.io_dataIn_2606(dataIn[2606]),
.io_dataIn_2607(dataIn[2607]),
.io_dataIn_2608(dataIn[2608]),
.io_dataIn_2609(dataIn[2609]),
.io_dataIn_2610(dataIn[2610]),
.io_dataIn_2611(dataIn[2611]),
.io_dataIn_2612(dataIn[2612]),
.io_dataIn_2613(dataIn[2613]),
.io_dataIn_2614(dataIn[2614]),
.io_dataIn_2615(dataIn[2615]),
.io_dataIn_2616(dataIn[2616]),
.io_dataIn_2617(dataIn[2617]),
.io_dataIn_2618(dataIn[2618]),
.io_dataIn_2619(dataIn[2619]),
.io_dataIn_2620(dataIn[2620]),
.io_dataIn_2621(dataIn[2621]),
.io_dataIn_2622(dataIn[2622]),
.io_dataIn_2623(dataIn[2623]),
.io_dataIn_2624(dataIn[2624]),
.io_dataIn_2625(dataIn[2625]),
.io_dataIn_2626(dataIn[2626]),
.io_dataIn_2627(dataIn[2627]),
.io_dataIn_2628(dataIn[2628]),
.io_dataIn_2629(dataIn[2629]),
.io_dataIn_2630(dataIn[2630]),
.io_dataIn_2631(dataIn[2631]),
.io_dataIn_2632(dataIn[2632]),
.io_dataIn_2633(dataIn[2633]),
.io_dataIn_2634(dataIn[2634]),
.io_dataIn_2635(dataIn[2635]),
.io_dataIn_2636(dataIn[2636]),
.io_dataIn_2637(dataIn[2637]),
.io_dataIn_2638(dataIn[2638]),
.io_dataIn_2639(dataIn[2639]),
.io_dataIn_2640(dataIn[2640]),
.io_dataIn_2641(dataIn[2641]),
.io_dataIn_2642(dataIn[2642]),
.io_dataIn_2643(dataIn[2643]),
.io_dataIn_2644(dataIn[2644]),
.io_dataIn_2645(dataIn[2645]),
.io_dataIn_2646(dataIn[2646]),
.io_dataIn_2647(dataIn[2647]),
.io_dataIn_2648(dataIn[2648]),
.io_dataIn_2649(dataIn[2649]),
.io_dataIn_2650(dataIn[2650]),
.io_dataIn_2651(dataIn[2651]),
.io_dataIn_2652(dataIn[2652]),
.io_dataIn_2653(dataIn[2653]),
.io_dataIn_2654(dataIn[2654]),
.io_dataIn_2655(dataIn[2655]),
.io_dataIn_2656(dataIn[2656]),
.io_dataIn_2657(dataIn[2657]),
.io_dataIn_2658(dataIn[2658]),
.io_dataIn_2659(dataIn[2659]),
.io_dataIn_2660(dataIn[2660]),
.io_dataIn_2661(dataIn[2661]),
.io_dataIn_2662(dataIn[2662]),
.io_dataIn_2663(dataIn[2663]),
.io_dataIn_2664(dataIn[2664]),
.io_dataIn_2665(dataIn[2665]),
.io_dataIn_2666(dataIn[2666]),
.io_dataIn_2667(dataIn[2667]),
.io_dataIn_2668(dataIn[2668]),
.io_dataIn_2669(dataIn[2669]),
.io_dataIn_2670(dataIn[2670]),
.io_dataIn_2671(dataIn[2671]),
.io_dataIn_2672(dataIn[2672]),
.io_dataIn_2673(dataIn[2673]),
.io_dataIn_2674(dataIn[2674]),
.io_dataIn_2675(dataIn[2675]),
.io_dataIn_2676(dataIn[2676]),
.io_dataIn_2677(dataIn[2677]),
.io_dataIn_2678(dataIn[2678]),
.io_dataIn_2679(dataIn[2679]),
.io_dataIn_2680(dataIn[2680]),
.io_dataIn_2681(dataIn[2681]),
.io_dataIn_2682(dataIn[2682]),
.io_dataIn_2683(dataIn[2683]),
.io_dataIn_2684(dataIn[2684]),
.io_dataIn_2685(dataIn[2685]),
.io_dataIn_2686(dataIn[2686]),
.io_dataIn_2687(dataIn[2687]),
.io_dataIn_2688(dataIn[2688]),
.io_dataIn_2689(dataIn[2689]),
.io_dataIn_2690(dataIn[2690]),
.io_dataIn_2691(dataIn[2691]),
.io_dataIn_2692(dataIn[2692]),
.io_dataIn_2693(dataIn[2693]),
.io_dataIn_2694(dataIn[2694]),
.io_dataIn_2695(dataIn[2695]),
.io_dataIn_2696(dataIn[2696]),
.io_dataIn_2697(dataIn[2697]),
.io_dataIn_2698(dataIn[2698]),
.io_dataIn_2699(dataIn[2699]),
.io_dataIn_2700(dataIn[2700]),
.io_dataIn_2701(dataIn[2701]),
.io_dataIn_2702(dataIn[2702]),
.io_dataIn_2703(dataIn[2703]),
.io_dataIn_2704(dataIn[2704]),
.io_dataIn_2705(dataIn[2705]),
.io_dataIn_2706(dataIn[2706]),
.io_dataIn_2707(dataIn[2707]),
.io_dataIn_2708(dataIn[2708]),
.io_dataIn_2709(dataIn[2709]),
.io_dataIn_2710(dataIn[2710]),
.io_dataIn_2711(dataIn[2711]),
.io_dataIn_2712(dataIn[2712]),
.io_dataIn_2713(dataIn[2713]),
.io_dataIn_2714(dataIn[2714]),
.io_dataIn_2715(dataIn[2715]),
.io_dataIn_2716(dataIn[2716]),
.io_dataIn_2717(dataIn[2717]),
.io_dataIn_2718(dataIn[2718]),
.io_dataIn_2719(dataIn[2719]),
.io_dataIn_2720(dataIn[2720]),
.io_dataIn_2721(dataIn[2721]),
.io_dataIn_2722(dataIn[2722]),
.io_dataIn_2723(dataIn[2723]),
.io_dataIn_2724(dataIn[2724]),
.io_dataIn_2725(dataIn[2725]),
.io_dataIn_2726(dataIn[2726]),
.io_dataIn_2727(dataIn[2727]),
.io_dataIn_2728(dataIn[2728]),
.io_dataIn_2729(dataIn[2729]),
.io_dataIn_2730(dataIn[2730]),
.io_dataIn_2731(dataIn[2731]),
.io_dataIn_2732(dataIn[2732]),
.io_dataIn_2733(dataIn[2733]),
.io_dataIn_2734(dataIn[2734]),
.io_dataIn_2735(dataIn[2735]),
.io_dataIn_2736(dataIn[2736]),
.io_dataIn_2737(dataIn[2737]),
.io_dataIn_2738(dataIn[2738]),
.io_dataIn_2739(dataIn[2739]),
.io_dataIn_2740(dataIn[2740]),
.io_dataIn_2741(dataIn[2741]),
.io_dataIn_2742(dataIn[2742]),
.io_dataIn_2743(dataIn[2743]),
.io_dataIn_2744(dataIn[2744]),
.io_dataIn_2745(dataIn[2745]),
.io_dataIn_2746(dataIn[2746]),
.io_dataIn_2747(dataIn[2747]),
.io_dataIn_2748(dataIn[2748]),
.io_dataIn_2749(dataIn[2749]),
.io_dataIn_2750(dataIn[2750]),
.io_dataIn_2751(dataIn[2751]),
.io_dataIn_2752(dataIn[2752]),
.io_dataIn_2753(dataIn[2753]),
.io_dataIn_2754(dataIn[2754]),
.io_dataIn_2755(dataIn[2755]),
.io_dataIn_2756(dataIn[2756]),
.io_dataIn_2757(dataIn[2757]),
.io_dataIn_2758(dataIn[2758]),
.io_dataIn_2759(dataIn[2759]),
.io_dataIn_2760(dataIn[2760]),
.io_dataIn_2761(dataIn[2761]),
.io_dataIn_2762(dataIn[2762]),
.io_dataIn_2763(dataIn[2763]),
.io_dataIn_2764(dataIn[2764]),
.io_dataIn_2765(dataIn[2765]),
.io_dataIn_2766(dataIn[2766]),
.io_dataIn_2767(dataIn[2767]),
.io_dataIn_2768(dataIn[2768]),
.io_dataIn_2769(dataIn[2769]),
.io_dataIn_2770(dataIn[2770]),
.io_dataIn_2771(dataIn[2771]),
.io_dataIn_2772(dataIn[2772]),
.io_dataIn_2773(dataIn[2773]),
.io_dataIn_2774(dataIn[2774]),
.io_dataIn_2775(dataIn[2775]),
.io_dataIn_2776(dataIn[2776]),
.io_dataIn_2777(dataIn[2777]),
.io_dataIn_2778(dataIn[2778]),
.io_dataIn_2779(dataIn[2779]),
.io_dataIn_2780(dataIn[2780]),
.io_dataIn_2781(dataIn[2781]),
.io_dataIn_2782(dataIn[2782]),
.io_dataIn_2783(dataIn[2783]),
.io_dataIn_2784(dataIn[2784]),
.io_dataIn_2785(dataIn[2785]),
.io_dataIn_2786(dataIn[2786]),
.io_dataIn_2787(dataIn[2787]),
.io_dataIn_2788(dataIn[2788]),
.io_dataIn_2789(dataIn[2789]),
.io_dataIn_2790(dataIn[2790]),
.io_dataIn_2791(dataIn[2791]),
.io_dataIn_2792(dataIn[2792]),
.io_dataIn_2793(dataIn[2793]),
.io_dataIn_2794(dataIn[2794]),
.io_dataIn_2795(dataIn[2795]),
.io_dataIn_2796(dataIn[2796]),
.io_dataIn_2797(dataIn[2797]),
.io_dataIn_2798(dataIn[2798]),
.io_dataIn_2799(dataIn[2799]),
.io_dataIn_2800(dataIn[2800]),
.io_dataIn_2801(dataIn[2801]),
.io_dataIn_2802(dataIn[2802]),
.io_dataIn_2803(dataIn[2803]),
.io_dataIn_2804(dataIn[2804]),
.io_dataIn_2805(dataIn[2805]),
.io_dataIn_2806(dataIn[2806]),
.io_dataIn_2807(dataIn[2807]),
.io_dataIn_2808(dataIn[2808]),
.io_dataIn_2809(dataIn[2809]),
.io_dataIn_2810(dataIn[2810]),
.io_dataIn_2811(dataIn[2811]),
.io_dataIn_2812(dataIn[2812]),
.io_dataIn_2813(dataIn[2813]),
.io_dataIn_2814(dataIn[2814]),
.io_dataIn_2815(dataIn[2815]),
.io_dataIn_2816(dataIn[2816]),
.io_dataIn_2817(dataIn[2817]),
.io_dataIn_2818(dataIn[2818]),
.io_dataIn_2819(dataIn[2819]),
.io_dataIn_2820(dataIn[2820]),
.io_dataIn_2821(dataIn[2821]),
.io_dataIn_2822(dataIn[2822]),
.io_dataIn_2823(dataIn[2823]),
.io_dataIn_2824(dataIn[2824]),
.io_dataIn_2825(dataIn[2825]),
.io_dataIn_2826(dataIn[2826]),
.io_dataIn_2827(dataIn[2827]),
.io_dataIn_2828(dataIn[2828]),
.io_dataIn_2829(dataIn[2829]),
.io_dataIn_2830(dataIn[2830]),
.io_dataIn_2831(dataIn[2831]),
.io_dataIn_2832(dataIn[2832]),
.io_dataIn_2833(dataIn[2833]),
.io_dataIn_2834(dataIn[2834]),
.io_dataIn_2835(dataIn[2835]),
.io_dataIn_2836(dataIn[2836]),
.io_dataIn_2837(dataIn[2837]),
.io_dataIn_2838(dataIn[2838]),
.io_dataIn_2839(dataIn[2839]),
.io_dataIn_2840(dataIn[2840]),
.io_dataIn_2841(dataIn[2841]),
.io_dataIn_2842(dataIn[2842]),
.io_dataIn_2843(dataIn[2843]),
.io_dataIn_2844(dataIn[2844]),
.io_dataIn_2845(dataIn[2845]),
.io_dataIn_2846(dataIn[2846]),
.io_dataIn_2847(dataIn[2847]),
.io_dataIn_2848(dataIn[2848]),
.io_dataIn_2849(dataIn[2849]),
.io_dataIn_2850(dataIn[2850]),
.io_dataIn_2851(dataIn[2851]),
.io_dataIn_2852(dataIn[2852]),
.io_dataIn_2853(dataIn[2853]),
.io_dataIn_2854(dataIn[2854]),
.io_dataIn_2855(dataIn[2855]),
.io_dataIn_2856(dataIn[2856]),
.io_dataIn_2857(dataIn[2857]),
.io_dataIn_2858(dataIn[2858]),
.io_dataIn_2859(dataIn[2859]),
.io_dataIn_2860(dataIn[2860]),
.io_dataIn_2861(dataIn[2861]),
.io_dataIn_2862(dataIn[2862]),
.io_dataIn_2863(dataIn[2863]),
.io_dataIn_2864(dataIn[2864]),
.io_dataIn_2865(dataIn[2865]),
.io_dataIn_2866(dataIn[2866]),
.io_dataIn_2867(dataIn[2867]),
.io_dataIn_2868(dataIn[2868]),
.io_dataIn_2869(dataIn[2869]),
.io_dataIn_2870(dataIn[2870]),
.io_dataIn_2871(dataIn[2871]),
.io_dataIn_2872(dataIn[2872]),
.io_dataIn_2873(dataIn[2873]),
.io_dataIn_2874(dataIn[2874]),
.io_dataIn_2875(dataIn[2875]),
.io_dataIn_2876(dataIn[2876]),
.io_dataIn_2877(dataIn[2877]),
.io_dataIn_2878(dataIn[2878]),
.io_dataIn_2879(dataIn[2879]),
.io_dataIn_2880(dataIn[2880]),
.io_dataIn_2881(dataIn[2881]),
.io_dataIn_2882(dataIn[2882]),
.io_dataIn_2883(dataIn[2883]),
.io_dataIn_2884(dataIn[2884]),
.io_dataIn_2885(dataIn[2885]),
.io_dataIn_2886(dataIn[2886]),
.io_dataIn_2887(dataIn[2887]),
.io_dataIn_2888(dataIn[2888]),
.io_dataIn_2889(dataIn[2889]),
.io_dataIn_2890(dataIn[2890]),
.io_dataIn_2891(dataIn[2891]),
.io_dataIn_2892(dataIn[2892]),
.io_dataIn_2893(dataIn[2893]),
.io_dataIn_2894(dataIn[2894]),
.io_dataIn_2895(dataIn[2895]),
.io_dataIn_2896(dataIn[2896]),
.io_dataIn_2897(dataIn[2897]),
.io_dataIn_2898(dataIn[2898]),
.io_dataIn_2899(dataIn[2899]),
.io_dataIn_2900(dataIn[2900]),
.io_dataIn_2901(dataIn[2901]),
.io_dataIn_2902(dataIn[2902]),
.io_dataIn_2903(dataIn[2903]),
.io_dataIn_2904(dataIn[2904]),
.io_dataIn_2905(dataIn[2905]),
.io_dataIn_2906(dataIn[2906]),
.io_dataIn_2907(dataIn[2907]),
.io_dataIn_2908(dataIn[2908]),
.io_dataIn_2909(dataIn[2909]),
.io_dataIn_2910(dataIn[2910]),
.io_dataIn_2911(dataIn[2911]),
.io_dataIn_2912(dataIn[2912]),
.io_dataIn_2913(dataIn[2913]),
.io_dataIn_2914(dataIn[2914]),
.io_dataIn_2915(dataIn[2915]),
.io_dataIn_2916(dataIn[2916]),
.io_dataIn_2917(dataIn[2917]),
.io_dataIn_2918(dataIn[2918]),
.io_dataIn_2919(dataIn[2919]),
.io_dataIn_2920(dataIn[2920]),
.io_dataIn_2921(dataIn[2921]),
.io_dataIn_2922(dataIn[2922]),
.io_dataIn_2923(dataIn[2923]),
.io_dataIn_2924(dataIn[2924]),
.io_dataIn_2925(dataIn[2925]),
.io_dataIn_2926(dataIn[2926]),
.io_dataIn_2927(dataIn[2927]),
.io_dataIn_2928(dataIn[2928]),
.io_dataIn_2929(dataIn[2929]),
.io_dataIn_2930(dataIn[2930]),
.io_dataIn_2931(dataIn[2931]),
.io_dataIn_2932(dataIn[2932]),
.io_dataIn_2933(dataIn[2933]),
.io_dataIn_2934(dataIn[2934]),
.io_dataIn_2935(dataIn[2935]),
.io_dataIn_2936(dataIn[2936]),
.io_dataIn_2937(dataIn[2937]),
.io_dataIn_2938(dataIn[2938]),
.io_dataIn_2939(dataIn[2939]),
.io_dataIn_2940(dataIn[2940]),
.io_dataIn_2941(dataIn[2941]),
.io_dataIn_2942(dataIn[2942]),
.io_dataIn_2943(dataIn[2943]),
.io_dataIn_2944(dataIn[2944]),
.io_dataIn_2945(dataIn[2945]),
.io_dataIn_2946(dataIn[2946]),
.io_dataIn_2947(dataIn[2947]),
.io_dataIn_2948(dataIn[2948]),
.io_dataIn_2949(dataIn[2949]),
.io_dataIn_2950(dataIn[2950]),
.io_dataIn_2951(dataIn[2951]),
.io_dataIn_2952(dataIn[2952]),
.io_dataIn_2953(dataIn[2953]),
.io_dataIn_2954(dataIn[2954]),
.io_dataIn_2955(dataIn[2955]),
.io_dataIn_2956(dataIn[2956]),
.io_dataIn_2957(dataIn[2957]),
.io_dataIn_2958(dataIn[2958]),
.io_dataIn_2959(dataIn[2959]),
.io_dataIn_2960(dataIn[2960]),
.io_dataIn_2961(dataIn[2961]),
.io_dataIn_2962(dataIn[2962]),
.io_dataIn_2963(dataIn[2963]),
.io_dataIn_2964(dataIn[2964]),
.io_dataIn_2965(dataIn[2965]),
.io_dataIn_2966(dataIn[2966]),
.io_dataIn_2967(dataIn[2967]),
.io_dataIn_2968(dataIn[2968]),
.io_dataIn_2969(dataIn[2969]),
.io_dataIn_2970(dataIn[2970]),
.io_dataIn_2971(dataIn[2971]),
.io_dataIn_2972(dataIn[2972]),
.io_dataIn_2973(dataIn[2973]),
.io_dataIn_2974(dataIn[2974]),
.io_dataIn_2975(dataIn[2975]),
.io_dataIn_2976(dataIn[2976]),
.io_dataIn_2977(dataIn[2977]),
.io_dataIn_2978(dataIn[2978]),
.io_dataIn_2979(dataIn[2979]),
.io_dataIn_2980(dataIn[2980]),
.io_dataIn_2981(dataIn[2981]),
.io_dataIn_2982(dataIn[2982]),
.io_dataIn_2983(dataIn[2983]),
.io_dataIn_2984(dataIn[2984]),
.io_dataIn_2985(dataIn[2985]),
.io_dataIn_2986(dataIn[2986]),
.io_dataIn_2987(dataIn[2987]),
.io_dataIn_2988(dataIn[2988]),
.io_dataIn_2989(dataIn[2989]),
.io_dataIn_2990(dataIn[2990]),
.io_dataIn_2991(dataIn[2991]),
.io_dataIn_2992(dataIn[2992]),
.io_dataIn_2993(dataIn[2993]),
.io_dataIn_2994(dataIn[2994]),
.io_dataIn_2995(dataIn[2995]),
.io_dataIn_2996(dataIn[2996]),
.io_dataIn_2997(dataIn[2997]),
.io_dataIn_2998(dataIn[2998]),
.io_dataIn_2999(dataIn[2999]),
.io_dataIn_3000(dataIn[3000]),
.io_dataIn_3001(dataIn[3001]),
.io_dataIn_3002(dataIn[3002]),
.io_dataIn_3003(dataIn[3003]),
.io_dataIn_3004(dataIn[3004]),
.io_dataIn_3005(dataIn[3005]),
.io_dataIn_3006(dataIn[3006]),
.io_dataIn_3007(dataIn[3007]),
.io_dataIn_3008(dataIn[3008]),
.io_dataIn_3009(dataIn[3009]),
.io_dataIn_3010(dataIn[3010]),
.io_dataIn_3011(dataIn[3011]),
.io_dataIn_3012(dataIn[3012]),
.io_dataIn_3013(dataIn[3013]),
.io_dataIn_3014(dataIn[3014]),
.io_dataIn_3015(dataIn[3015]),
.io_dataIn_3016(dataIn[3016]),
.io_dataIn_3017(dataIn[3017]),
.io_dataIn_3018(dataIn[3018]),
.io_dataIn_3019(dataIn[3019]),
.io_dataIn_3020(dataIn[3020]),
.io_dataIn_3021(dataIn[3021]),
.io_dataIn_3022(dataIn[3022]),
.io_dataIn_3023(dataIn[3023]),
.io_dataIn_3024(dataIn[3024]),
.io_dataIn_3025(dataIn[3025]),
.io_dataIn_3026(dataIn[3026]),
.io_dataIn_3027(dataIn[3027]),
.io_dataIn_3028(dataIn[3028]),
.io_dataIn_3029(dataIn[3029]),
.io_dataIn_3030(dataIn[3030]),
.io_dataIn_3031(dataIn[3031]),
.io_dataIn_3032(dataIn[3032]),
.io_dataIn_3033(dataIn[3033]),
.io_dataIn_3034(dataIn[3034]),
.io_dataIn_3035(dataIn[3035]),
.io_dataIn_3036(dataIn[3036]),
.io_dataIn_3037(dataIn[3037]),
.io_dataIn_3038(dataIn[3038]),
.io_dataIn_3039(dataIn[3039]),
.io_dataIn_3040(dataIn[3040]),
.io_dataIn_3041(dataIn[3041]),
.io_dataIn_3042(dataIn[3042]),
.io_dataIn_3043(dataIn[3043]),
.io_dataIn_3044(dataIn[3044]),
.io_dataIn_3045(dataIn[3045]),
.io_dataIn_3046(dataIn[3046]),
.io_dataIn_3047(dataIn[3047]),
.io_dataIn_3048(dataIn[3048]),
.io_dataIn_3049(dataIn[3049]),
.io_dataIn_3050(dataIn[3050]),
.io_dataIn_3051(dataIn[3051]),
.io_dataIn_3052(dataIn[3052]),
.io_dataIn_3053(dataIn[3053]),
.io_dataIn_3054(dataIn[3054]),
.io_dataIn_3055(dataIn[3055]),
.io_dataIn_3056(dataIn[3056]),
.io_dataIn_3057(dataIn[3057]),
.io_dataIn_3058(dataIn[3058]),
.io_dataIn_3059(dataIn[3059]),
.io_dataIn_3060(dataIn[3060]),
.io_dataIn_3061(dataIn[3061]),
.io_dataIn_3062(dataIn[3062]),
.io_dataIn_3063(dataIn[3063]),
.io_dataIn_3064(dataIn[3064]),
.io_dataIn_3065(dataIn[3065]),
.io_dataIn_3066(dataIn[3066]),
.io_dataIn_3067(dataIn[3067]),
.io_dataIn_3068(dataIn[3068]),
.io_dataIn_3069(dataIn[3069]),
.io_dataIn_3070(dataIn[3070]),
.io_dataIn_3071(dataIn[3071]),
.io_dataIn_3072(dataIn[3072]),
.io_dataIn_3073(dataIn[3073]),
.io_dataIn_3074(dataIn[3074]),
.io_dataIn_3075(dataIn[3075]),
.io_dataIn_3076(dataIn[3076]),
.io_dataIn_3077(dataIn[3077]),
.io_dataIn_3078(dataIn[3078]),
.io_dataIn_3079(dataIn[3079]),
.io_dataIn_3080(dataIn[3080]),
.io_dataIn_3081(dataIn[3081]),
.io_dataIn_3082(dataIn[3082]),
.io_dataIn_3083(dataIn[3083]),
.io_dataIn_3084(dataIn[3084]),
.io_dataIn_3085(dataIn[3085]),
.io_dataIn_3086(dataIn[3086]),
.io_dataIn_3087(dataIn[3087]),
.io_dataIn_3088(dataIn[3088]),
.io_dataIn_3089(dataIn[3089]),
.io_dataIn_3090(dataIn[3090]),
.io_dataIn_3091(dataIn[3091]),
.io_dataIn_3092(dataIn[3092]),
.io_dataIn_3093(dataIn[3093]),
.io_dataIn_3094(dataIn[3094]),
.io_dataIn_3095(dataIn[3095]),
.io_dataIn_3096(dataIn[3096]),
.io_dataIn_3097(dataIn[3097]),
.io_dataIn_3098(dataIn[3098]),
.io_dataIn_3099(dataIn[3099]),
.io_dataIn_3100(dataIn[3100]),
.io_dataIn_3101(dataIn[3101]),
.io_dataIn_3102(dataIn[3102]),
.io_dataIn_3103(dataIn[3103]),
.io_dataIn_3104(dataIn[3104]),
.io_dataIn_3105(dataIn[3105]),
.io_dataIn_3106(dataIn[3106]),
.io_dataIn_3107(dataIn[3107]),
.io_dataIn_3108(dataIn[3108]),
.io_dataIn_3109(dataIn[3109]),
.io_dataIn_3110(dataIn[3110]),
.io_dataIn_3111(dataIn[3111]),
.io_dataIn_3112(dataIn[3112]),
.io_dataIn_3113(dataIn[3113]),
.io_dataIn_3114(dataIn[3114]),
.io_dataIn_3115(dataIn[3115]),
.io_dataIn_3116(dataIn[3116]),
.io_dataIn_3117(dataIn[3117]),
.io_dataIn_3118(dataIn[3118]),
.io_dataIn_3119(dataIn[3119]),
.io_dataIn_3120(dataIn[3120]),
.io_dataIn_3121(dataIn[3121]),
.io_dataIn_3122(dataIn[3122]),
.io_dataIn_3123(dataIn[3123]),
.io_dataIn_3124(dataIn[3124]),
.io_dataIn_3125(dataIn[3125]),
.io_dataIn_3126(dataIn[3126]),
.io_dataIn_3127(dataIn[3127]),
.io_dataIn_3128(dataIn[3128]),
.io_dataIn_3129(dataIn[3129]),
.io_dataIn_3130(dataIn[3130]),
.io_dataIn_3131(dataIn[3131]),
.io_dataIn_3132(dataIn[3132]),
.io_dataIn_3133(dataIn[3133]),
.io_dataIn_3134(dataIn[3134]),
.io_dataIn_3135(dataIn[3135]),
.io_dataIn_3136(dataIn[3136]),
.io_dataIn_3137(dataIn[3137]),
.io_dataIn_3138(dataIn[3138]),
.io_dataIn_3139(dataIn[3139]),
.io_dataIn_3140(dataIn[3140]),
.io_dataIn_3141(dataIn[3141]),
.io_dataIn_3142(dataIn[3142]),
.io_dataIn_3143(dataIn[3143]),
.io_dataIn_3144(dataIn[3144]),
.io_dataIn_3145(dataIn[3145]),
.io_dataIn_3146(dataIn[3146]),
.io_dataIn_3147(dataIn[3147]),
.io_dataIn_3148(dataIn[3148]),
.io_dataIn_3149(dataIn[3149]),
.io_dataIn_3150(dataIn[3150]),
.io_dataIn_3151(dataIn[3151]),
.io_dataIn_3152(dataIn[3152]),
.io_dataIn_3153(dataIn[3153]),
.io_dataIn_3154(dataIn[3154]),
.io_dataIn_3155(dataIn[3155]),
.io_dataIn_3156(dataIn[3156]),
.io_dataIn_3157(dataIn[3157]),
.io_dataIn_3158(dataIn[3158]),
.io_dataIn_3159(dataIn[3159]),
.io_dataIn_3160(dataIn[3160]),
.io_dataIn_3161(dataIn[3161]),
.io_dataIn_3162(dataIn[3162]),
.io_dataIn_3163(dataIn[3163]),
.io_dataIn_3164(dataIn[3164]),
.io_dataIn_3165(dataIn[3165]),
.io_dataIn_3166(dataIn[3166]),
.io_dataIn_3167(dataIn[3167]),
.io_dataIn_3168(dataIn[3168]),
.io_dataIn_3169(dataIn[3169]),
.io_dataIn_3170(dataIn[3170]),
.io_dataIn_3171(dataIn[3171]),
.io_dataIn_3172(dataIn[3172]),
.io_dataIn_3173(dataIn[3173]),
.io_dataIn_3174(dataIn[3174]),
.io_dataIn_3175(dataIn[3175]),
.io_dataIn_3176(dataIn[3176]),
.io_dataIn_3177(dataIn[3177]),
.io_dataIn_3178(dataIn[3178]),
.io_dataIn_3179(dataIn[3179]),
.io_dataIn_3180(dataIn[3180]),
.io_dataIn_3181(dataIn[3181]),
.io_dataIn_3182(dataIn[3182]),
.io_dataIn_3183(dataIn[3183]),
.io_dataIn_3184(dataIn[3184]),
.io_dataIn_3185(dataIn[3185]),
.io_dataIn_3186(dataIn[3186]),
.io_dataIn_3187(dataIn[3187]),
.io_dataIn_3188(dataIn[3188]),
.io_dataIn_3189(dataIn[3189]),
.io_dataIn_3190(dataIn[3190]),
.io_dataIn_3191(dataIn[3191]),
.io_dataIn_3192(dataIn[3192]),
.io_dataIn_3193(dataIn[3193]),
.io_dataIn_3194(dataIn[3194]),
.io_dataIn_3195(dataIn[3195]),
.io_dataIn_3196(dataIn[3196]),
.io_dataIn_3197(dataIn[3197]),
.io_dataIn_3198(dataIn[3198]),
.io_dataIn_3199(dataIn[3199]),
.io_dataIn_3200(dataIn[3200]),
.io_dataIn_3201(dataIn[3201]),
.io_dataIn_3202(dataIn[3202]),
.io_dataIn_3203(dataIn[3203]),
.io_dataIn_3204(dataIn[3204]),
.io_dataIn_3205(dataIn[3205]),
.io_dataIn_3206(dataIn[3206]),
.io_dataIn_3207(dataIn[3207]),
.io_dataIn_3208(dataIn[3208]),
.io_dataIn_3209(dataIn[3209]),
.io_dataIn_3210(dataIn[3210]),
.io_dataIn_3211(dataIn[3211]),
.io_dataIn_3212(dataIn[3212]),
.io_dataIn_3213(dataIn[3213]),
.io_dataIn_3214(dataIn[3214]),
.io_dataIn_3215(dataIn[3215]),
.io_dataIn_3216(dataIn[3216]),
.io_dataIn_3217(dataIn[3217]),
.io_dataIn_3218(dataIn[3218]),
.io_dataIn_3219(dataIn[3219]),
.io_dataIn_3220(dataIn[3220]),
.io_dataIn_3221(dataIn[3221]),
.io_dataIn_3222(dataIn[3222]),
.io_dataIn_3223(dataIn[3223]),
.io_dataIn_3224(dataIn[3224]),
.io_dataIn_3225(dataIn[3225]),
.io_dataIn_3226(dataIn[3226]),
.io_dataIn_3227(dataIn[3227]),
.io_dataIn_3228(dataIn[3228]),
.io_dataIn_3229(dataIn[3229]),
.io_dataIn_3230(dataIn[3230]),
.io_dataIn_3231(dataIn[3231]),
.io_dataIn_3232(dataIn[3232]),
.io_dataIn_3233(dataIn[3233]),
.io_dataIn_3234(dataIn[3234]),
.io_dataIn_3235(dataIn[3235]),
.io_dataIn_3236(dataIn[3236]),
.io_dataIn_3237(dataIn[3237]),
.io_dataIn_3238(dataIn[3238]),
.io_dataIn_3239(dataIn[3239]),
.io_dataIn_3240(dataIn[3240]),
.io_dataIn_3241(dataIn[3241]),
.io_dataIn_3242(dataIn[3242]),
.io_dataIn_3243(dataIn[3243]),
.io_dataIn_3244(dataIn[3244]),
.io_dataIn_3245(dataIn[3245]),
.io_dataIn_3246(dataIn[3246]),
.io_dataIn_3247(dataIn[3247]),
.io_dataIn_3248(dataIn[3248]),
.io_dataIn_3249(dataIn[3249]),
.io_dataIn_3250(dataIn[3250]),
.io_dataIn_3251(dataIn[3251]),
.io_dataIn_3252(dataIn[3252]),
.io_dataIn_3253(dataIn[3253]),
.io_dataIn_3254(dataIn[3254]),
.io_dataIn_3255(dataIn[3255]),
.io_dataIn_3256(dataIn[3256]),
.io_dataIn_3257(dataIn[3257]),
.io_dataIn_3258(dataIn[3258]),
.io_dataIn_3259(dataIn[3259]),
.io_dataIn_3260(dataIn[3260]),
.io_dataIn_3261(dataIn[3261]),
.io_dataIn_3262(dataIn[3262]),
.io_dataIn_3263(dataIn[3263]),
.io_dataIn_3264(dataIn[3264]),
.io_dataIn_3265(dataIn[3265]),
.io_dataIn_3266(dataIn[3266]),
.io_dataIn_3267(dataIn[3267]),
.io_dataIn_3268(dataIn[3268]),
.io_dataIn_3269(dataIn[3269]),
.io_dataIn_3270(dataIn[3270]),
.io_dataIn_3271(dataIn[3271]),
.io_dataIn_3272(dataIn[3272]),
.io_dataIn_3273(dataIn[3273]),
.io_dataIn_3274(dataIn[3274]),
.io_dataIn_3275(dataIn[3275]),
.io_dataIn_3276(dataIn[3276]),
.io_dataIn_3277(dataIn[3277]),
.io_dataIn_3278(dataIn[3278]),
.io_dataIn_3279(dataIn[3279]),
.io_dataIn_3280(dataIn[3280]),
.io_dataIn_3281(dataIn[3281]),
.io_dataIn_3282(dataIn[3282]),
.io_dataIn_3283(dataIn[3283]),
.io_dataIn_3284(dataIn[3284]),
.io_dataIn_3285(dataIn[3285]),
.io_dataIn_3286(dataIn[3286]),
.io_dataIn_3287(dataIn[3287]),
.io_dataIn_3288(dataIn[3288]),
.io_dataIn_3289(dataIn[3289]),
.io_dataIn_3290(dataIn[3290]),
.io_dataIn_3291(dataIn[3291]),
.io_dataIn_3292(dataIn[3292]),
.io_dataIn_3293(dataIn[3293]),
.io_dataIn_3294(dataIn[3294]),
.io_dataIn_3295(dataIn[3295]),
.io_dataIn_3296(dataIn[3296]),
.io_dataIn_3297(dataIn[3297]),
.io_dataIn_3298(dataIn[3298]),
.io_dataIn_3299(dataIn[3299]),
.io_dataIn_3300(dataIn[3300]),
.io_dataIn_3301(dataIn[3301]),
.io_dataIn_3302(dataIn[3302]),
.io_dataIn_3303(dataIn[3303]),
.io_dataIn_3304(dataIn[3304]),
.io_dataIn_3305(dataIn[3305]),
.io_dataIn_3306(dataIn[3306]),
.io_dataIn_3307(dataIn[3307]),
.io_dataIn_3308(dataIn[3308]),
.io_dataIn_3309(dataIn[3309]),
.io_dataIn_3310(dataIn[3310]),
.io_dataIn_3311(dataIn[3311]),
.io_dataIn_3312(dataIn[3312]),
.io_dataIn_3313(dataIn[3313]),
.io_dataIn_3314(dataIn[3314]),
.io_dataIn_3315(dataIn[3315]),
.io_dataIn_3316(dataIn[3316]),
.io_dataIn_3317(dataIn[3317]),
.io_dataIn_3318(dataIn[3318]),
.io_dataIn_3319(dataIn[3319]),
.io_dataIn_3320(dataIn[3320]),
.io_dataIn_3321(dataIn[3321]),
.io_dataIn_3322(dataIn[3322]),
.io_dataIn_3323(dataIn[3323]),
.io_dataIn_3324(dataIn[3324]),
.io_dataIn_3325(dataIn[3325]),
.io_dataIn_3326(dataIn[3326]),
.io_dataIn_3327(dataIn[3327]),
.io_dataIn_3328(dataIn[3328]),
.io_dataIn_3329(dataIn[3329]),
.io_dataIn_3330(dataIn[3330]),
.io_dataIn_3331(dataIn[3331]),
.io_dataIn_3332(dataIn[3332]),
.io_dataIn_3333(dataIn[3333]),
.io_dataIn_3334(dataIn[3334]),
.io_dataIn_3335(dataIn[3335]),
.io_dataIn_3336(dataIn[3336]),
.io_dataIn_3337(dataIn[3337]),
.io_dataIn_3338(dataIn[3338]),
.io_dataIn_3339(dataIn[3339]),
.io_dataIn_3340(dataIn[3340]),
.io_dataIn_3341(dataIn[3341]),
.io_dataIn_3342(dataIn[3342]),
.io_dataIn_3343(dataIn[3343]),
.io_dataIn_3344(dataIn[3344]),
.io_dataIn_3345(dataIn[3345]),
.io_dataIn_3346(dataIn[3346]),
.io_dataIn_3347(dataIn[3347]),
.io_dataIn_3348(dataIn[3348]),
.io_dataIn_3349(dataIn[3349]),
.io_dataIn_3350(dataIn[3350]),
.io_dataIn_3351(dataIn[3351]),
.io_dataIn_3352(dataIn[3352]),
.io_dataIn_3353(dataIn[3353]),
.io_dataIn_3354(dataIn[3354]),
.io_dataIn_3355(dataIn[3355]),
.io_dataIn_3356(dataIn[3356]),
.io_dataIn_3357(dataIn[3357]),
.io_dataIn_3358(dataIn[3358]),
.io_dataIn_3359(dataIn[3359]),
.io_dataIn_3360(dataIn[3360]),
.io_dataIn_3361(dataIn[3361]),
.io_dataIn_3362(dataIn[3362]),
.io_dataIn_3363(dataIn[3363]),
.io_dataIn_3364(dataIn[3364]),
.io_dataIn_3365(dataIn[3365]),
.io_dataIn_3366(dataIn[3366]),
.io_dataIn_3367(dataIn[3367]),
.io_dataIn_3368(dataIn[3368]),
.io_dataIn_3369(dataIn[3369]),
.io_dataIn_3370(dataIn[3370]),
.io_dataIn_3371(dataIn[3371]),
.io_dataIn_3372(dataIn[3372]),
.io_dataIn_3373(dataIn[3373]),
.io_dataIn_3374(dataIn[3374]),
.io_dataIn_3375(dataIn[3375]),
.io_dataIn_3376(dataIn[3376]),
.io_dataIn_3377(dataIn[3377]),
.io_dataIn_3378(dataIn[3378]),
.io_dataIn_3379(dataIn[3379]),
.io_dataIn_3380(dataIn[3380]),
.io_dataIn_3381(dataIn[3381]),
.io_dataIn_3382(dataIn[3382]),
.io_dataIn_3383(dataIn[3383]),
.io_dataIn_3384(dataIn[3384]),
.io_dataIn_3385(dataIn[3385]),
.io_dataIn_3386(dataIn[3386]),
.io_dataIn_3387(dataIn[3387]),
.io_dataIn_3388(dataIn[3388]),
.io_dataIn_3389(dataIn[3389]),
.io_dataIn_3390(dataIn[3390]),
.io_dataIn_3391(dataIn[3391]),
.io_dataIn_3392(dataIn[3392]),
.io_dataIn_3393(dataIn[3393]),
.io_dataIn_3394(dataIn[3394]),
.io_dataIn_3395(dataIn[3395]),
.io_dataIn_3396(dataIn[3396]),
.io_dataIn_3397(dataIn[3397]),
.io_dataIn_3398(dataIn[3398]),
.io_dataIn_3399(dataIn[3399]),
.io_dataIn_3400(dataIn[3400]),
.io_dataIn_3401(dataIn[3401]),
.io_dataIn_3402(dataIn[3402]),
.io_dataIn_3403(dataIn[3403]),
.io_dataIn_3404(dataIn[3404]),
.io_dataIn_3405(dataIn[3405]),
.io_dataIn_3406(dataIn[3406]),
.io_dataIn_3407(dataIn[3407]),
.io_dataIn_3408(dataIn[3408]),
.io_dataIn_3409(dataIn[3409]),
.io_dataIn_3410(dataIn[3410]),
.io_dataIn_3411(dataIn[3411]),
.io_dataIn_3412(dataIn[3412]),
.io_dataIn_3413(dataIn[3413]),
.io_dataIn_3414(dataIn[3414]),
.io_dataIn_3415(dataIn[3415]),
.io_dataIn_3416(dataIn[3416]),
.io_dataIn_3417(dataIn[3417]),
.io_dataIn_3418(dataIn[3418]),
.io_dataIn_3419(dataIn[3419]),
.io_dataIn_3420(dataIn[3420]),
.io_dataIn_3421(dataIn[3421]),
.io_dataIn_3422(dataIn[3422]),
.io_dataIn_3423(dataIn[3423]),
.io_dataIn_3424(dataIn[3424]),
.io_dataIn_3425(dataIn[3425]),
.io_dataIn_3426(dataIn[3426]),
.io_dataIn_3427(dataIn[3427]),
.io_dataIn_3428(dataIn[3428]),
.io_dataIn_3429(dataIn[3429]),
.io_dataIn_3430(dataIn[3430]),
.io_dataIn_3431(dataIn[3431]),
.io_dataIn_3432(dataIn[3432]),
.io_dataIn_3433(dataIn[3433]),
.io_dataIn_3434(dataIn[3434]),
.io_dataIn_3435(dataIn[3435]),
.io_dataIn_3436(dataIn[3436]),
.io_dataIn_3437(dataIn[3437]),
.io_dataIn_3438(dataIn[3438]),
.io_dataIn_3439(dataIn[3439]),
.io_dataIn_3440(dataIn[3440]),
.io_dataIn_3441(dataIn[3441]),
.io_dataIn_3442(dataIn[3442]),
.io_dataIn_3443(dataIn[3443]),
.io_dataIn_3444(dataIn[3444]),
.io_dataIn_3445(dataIn[3445]),
.io_dataIn_3446(dataIn[3446]),
.io_dataIn_3447(dataIn[3447]),
.io_dataIn_3448(dataIn[3448]),
.io_dataIn_3449(dataIn[3449]),
.io_dataIn_3450(dataIn[3450]),
.io_dataIn_3451(dataIn[3451]),
.io_dataIn_3452(dataIn[3452]),
.io_dataIn_3453(dataIn[3453]),
.io_dataIn_3454(dataIn[3454]),
.io_dataIn_3455(dataIn[3455]),
.io_dataIn_3456(dataIn[3456]),
.io_dataIn_3457(dataIn[3457]),
.io_dataIn_3458(dataIn[3458]),
.io_dataIn_3459(dataIn[3459]),
.io_dataIn_3460(dataIn[3460]),
.io_dataIn_3461(dataIn[3461]),
.io_dataIn_3462(dataIn[3462]),
.io_dataIn_3463(dataIn[3463]),
.io_dataIn_3464(dataIn[3464]),
.io_dataIn_3465(dataIn[3465]),
.io_dataIn_3466(dataIn[3466]),
.io_dataIn_3467(dataIn[3467]),
.io_dataIn_3468(dataIn[3468]),
.io_dataIn_3469(dataIn[3469]),
.io_dataIn_3470(dataIn[3470]),
.io_dataIn_3471(dataIn[3471]),
.io_dataIn_3472(dataIn[3472]),
.io_dataIn_3473(dataIn[3473]),
.io_dataIn_3474(dataIn[3474]),
.io_dataIn_3475(dataIn[3475]),
.io_dataIn_3476(dataIn[3476]),
.io_dataIn_3477(dataIn[3477]),
.io_dataIn_3478(dataIn[3478]),
.io_dataIn_3479(dataIn[3479]),
.io_dataIn_3480(dataIn[3480]),
.io_dataIn_3481(dataIn[3481]),
.io_dataIn_3482(dataIn[3482]),
.io_dataIn_3483(dataIn[3483]),
.io_dataIn_3484(dataIn[3484]),
.io_dataIn_3485(dataIn[3485]),
.io_dataIn_3486(dataIn[3486]),
.io_dataIn_3487(dataIn[3487]),
.io_dataIn_3488(dataIn[3488]),
.io_dataIn_3489(dataIn[3489]),
.io_dataIn_3490(dataIn[3490]),
.io_dataIn_3491(dataIn[3491]),
.io_dataIn_3492(dataIn[3492]),
.io_dataIn_3493(dataIn[3493]),
.io_dataIn_3494(dataIn[3494]),
.io_dataIn_3495(dataIn[3495]),
.io_dataIn_3496(dataIn[3496]),
.io_dataIn_3497(dataIn[3497]),
.io_dataIn_3498(dataIn[3498]),
.io_dataIn_3499(dataIn[3499]),
.io_dataIn_3500(dataIn[3500]),
.io_dataIn_3501(dataIn[3501]),
.io_dataIn_3502(dataIn[3502]),
.io_dataIn_3503(dataIn[3503]),
.io_dataIn_3504(dataIn[3504]),
.io_dataIn_3505(dataIn[3505]),
.io_dataIn_3506(dataIn[3506]),
.io_dataIn_3507(dataIn[3507]),
.io_dataIn_3508(dataIn[3508]),
.io_dataIn_3509(dataIn[3509]),
.io_dataIn_3510(dataIn[3510]),
.io_dataIn_3511(dataIn[3511]),
.io_dataIn_3512(dataIn[3512]),
.io_dataIn_3513(dataIn[3513]),
.io_dataIn_3514(dataIn[3514]),
.io_dataIn_3515(dataIn[3515]),
.io_dataIn_3516(dataIn[3516]),
.io_dataIn_3517(dataIn[3517]),
.io_dataIn_3518(dataIn[3518]),
.io_dataIn_3519(dataIn[3519]),
.io_dataIn_3520(dataIn[3520]),
.io_dataIn_3521(dataIn[3521]),
.io_dataIn_3522(dataIn[3522]),
.io_dataIn_3523(dataIn[3523]),
.io_dataIn_3524(dataIn[3524]),
.io_dataIn_3525(dataIn[3525]),
.io_dataIn_3526(dataIn[3526]),
.io_dataIn_3527(dataIn[3527]),
.io_dataIn_3528(dataIn[3528]),
.io_dataIn_3529(dataIn[3529]),
.io_dataIn_3530(dataIn[3530]),
.io_dataIn_3531(dataIn[3531]),
.io_dataIn_3532(dataIn[3532]),
.io_dataIn_3533(dataIn[3533]),
.io_dataIn_3534(dataIn[3534]),
.io_dataIn_3535(dataIn[3535]),
.io_dataIn_3536(dataIn[3536]),
.io_dataIn_3537(dataIn[3537]),
.io_dataIn_3538(dataIn[3538]),
.io_dataIn_3539(dataIn[3539]),
.io_dataIn_3540(dataIn[3540]),
.io_dataIn_3541(dataIn[3541]),
.io_dataIn_3542(dataIn[3542]),
.io_dataIn_3543(dataIn[3543]),
.io_dataIn_3544(dataIn[3544]),
.io_dataIn_3545(dataIn[3545]),
.io_dataIn_3546(dataIn[3546]),
.io_dataIn_3547(dataIn[3547]),
.io_dataIn_3548(dataIn[3548]),
.io_dataIn_3549(dataIn[3549]),
.io_dataIn_3550(dataIn[3550]),
.io_dataIn_3551(dataIn[3551]),
.io_dataIn_3552(dataIn[3552]),
.io_dataIn_3553(dataIn[3553]),
.io_dataIn_3554(dataIn[3554]),
.io_dataIn_3555(dataIn[3555]),
.io_dataIn_3556(dataIn[3556]),
.io_dataIn_3557(dataIn[3557]),
.io_dataIn_3558(dataIn[3558]),
.io_dataIn_3559(dataIn[3559]),
.io_dataIn_3560(dataIn[3560]),
.io_dataIn_3561(dataIn[3561]),
.io_dataIn_3562(dataIn[3562]),
.io_dataIn_3563(dataIn[3563]),
.io_dataIn_3564(dataIn[3564]),
.io_dataIn_3565(dataIn[3565]),
.io_dataIn_3566(dataIn[3566]),
.io_dataIn_3567(dataIn[3567]),
.io_dataIn_3568(dataIn[3568]),
.io_dataIn_3569(dataIn[3569]),
.io_dataIn_3570(dataIn[3570]),
.io_dataIn_3571(dataIn[3571]),
.io_dataIn_3572(dataIn[3572]),
.io_dataIn_3573(dataIn[3573]),
.io_dataIn_3574(dataIn[3574]),
.io_dataIn_3575(dataIn[3575]),
.io_dataIn_3576(dataIn[3576]),
.io_dataIn_3577(dataIn[3577]),
.io_dataIn_3578(dataIn[3578]),
.io_dataIn_3579(dataIn[3579]),
.io_dataIn_3580(dataIn[3580]),
.io_dataIn_3581(dataIn[3581]),
.io_dataIn_3582(dataIn[3582]),
.io_dataIn_3583(dataIn[3583]),
.io_dataIn_3584(dataIn[3584]),
.io_dataIn_3585(dataIn[3585]),
.io_dataIn_3586(dataIn[3586]),
.io_dataIn_3587(dataIn[3587]),
.io_dataIn_3588(dataIn[3588]),
.io_dataIn_3589(dataIn[3589]),
.io_dataIn_3590(dataIn[3590]),
.io_dataIn_3591(dataIn[3591]),
.io_dataIn_3592(dataIn[3592]),
.io_dataIn_3593(dataIn[3593]),
.io_dataIn_3594(dataIn[3594]),
.io_dataIn_3595(dataIn[3595]),
.io_dataIn_3596(dataIn[3596]),
.io_dataIn_3597(dataIn[3597]),
.io_dataIn_3598(dataIn[3598]),
.io_dataIn_3599(dataIn[3599]),
.io_dataIn_3600(dataIn[3600]),
.io_dataIn_3601(dataIn[3601]),
.io_dataIn_3602(dataIn[3602]),
.io_dataIn_3603(dataIn[3603]),
.io_dataIn_3604(dataIn[3604]),
.io_dataIn_3605(dataIn[3605]),
.io_dataIn_3606(dataIn[3606]),
.io_dataIn_3607(dataIn[3607]),
.io_dataIn_3608(dataIn[3608]),
.io_dataIn_3609(dataIn[3609]),
.io_dataIn_3610(dataIn[3610]),
.io_dataIn_3611(dataIn[3611]),
.io_dataIn_3612(dataIn[3612]),
.io_dataIn_3613(dataIn[3613]),
.io_dataIn_3614(dataIn[3614]),
.io_dataIn_3615(dataIn[3615]),
.io_dataIn_3616(dataIn[3616]),
.io_dataIn_3617(dataIn[3617]),
.io_dataIn_3618(dataIn[3618]),
.io_dataIn_3619(dataIn[3619]),
.io_dataIn_3620(dataIn[3620]),
.io_dataIn_3621(dataIn[3621]),
.io_dataIn_3622(dataIn[3622]),
.io_dataIn_3623(dataIn[3623]),
.io_dataIn_3624(dataIn[3624]),
.io_dataIn_3625(dataIn[3625]),
.io_dataIn_3626(dataIn[3626]),
.io_dataIn_3627(dataIn[3627]),
.io_dataIn_3628(dataIn[3628]),
.io_dataIn_3629(dataIn[3629]),
.io_dataIn_3630(dataIn[3630]),
.io_dataIn_3631(dataIn[3631]),
.io_dataIn_3632(dataIn[3632]),
.io_dataIn_3633(dataIn[3633]),
.io_dataIn_3634(dataIn[3634]),
.io_dataIn_3635(dataIn[3635]),
.io_dataIn_3636(dataIn[3636]),
.io_dataIn_3637(dataIn[3637]),
.io_dataIn_3638(dataIn[3638]),
.io_dataIn_3639(dataIn[3639]),
.io_dataIn_3640(dataIn[3640]),
.io_dataIn_3641(dataIn[3641]),
.io_dataIn_3642(dataIn[3642]),
.io_dataIn_3643(dataIn[3643]),
.io_dataIn_3644(dataIn[3644]),
.io_dataIn_3645(dataIn[3645]),
.io_dataIn_3646(dataIn[3646]),
.io_dataIn_3647(dataIn[3647]),
.io_dataIn_3648(dataIn[3648]),
.io_dataIn_3649(dataIn[3649]),
.io_dataIn_3650(dataIn[3650]),
.io_dataIn_3651(dataIn[3651]),
.io_dataIn_3652(dataIn[3652]),
.io_dataIn_3653(dataIn[3653]),
.io_dataIn_3654(dataIn[3654]),
.io_dataIn_3655(dataIn[3655]),
.io_dataIn_3656(dataIn[3656]),
.io_dataIn_3657(dataIn[3657]),
.io_dataIn_3658(dataIn[3658]),
.io_dataIn_3659(dataIn[3659]),
.io_dataIn_3660(dataIn[3660]),
.io_dataIn_3661(dataIn[3661]),
.io_dataIn_3662(dataIn[3662]),
.io_dataIn_3663(dataIn[3663]),
.io_dataIn_3664(dataIn[3664]),
.io_dataIn_3665(dataIn[3665]),
.io_dataIn_3666(dataIn[3666]),
.io_dataIn_3667(dataIn[3667]),
.io_dataIn_3668(dataIn[3668]),
.io_dataIn_3669(dataIn[3669]),
.io_dataIn_3670(dataIn[3670]),
.io_dataIn_3671(dataIn[3671]),
.io_dataIn_3672(dataIn[3672]),
.io_dataIn_3673(dataIn[3673]),
.io_dataIn_3674(dataIn[3674]),
.io_dataIn_3675(dataIn[3675]),
.io_dataIn_3676(dataIn[3676]),
.io_dataIn_3677(dataIn[3677]),
.io_dataIn_3678(dataIn[3678]),
.io_dataIn_3679(dataIn[3679]),
.io_dataIn_3680(dataIn[3680]),
.io_dataIn_3681(dataIn[3681]),
.io_dataIn_3682(dataIn[3682]),
.io_dataIn_3683(dataIn[3683]),
.io_dataIn_3684(dataIn[3684]),
.io_dataIn_3685(dataIn[3685]),
.io_dataIn_3686(dataIn[3686]),
.io_dataIn_3687(dataIn[3687]),
.io_dataIn_3688(dataIn[3688]),
.io_dataIn_3689(dataIn[3689]),
.io_dataIn_3690(dataIn[3690]),
.io_dataIn_3691(dataIn[3691]),
.io_dataIn_3692(dataIn[3692]),
.io_dataIn_3693(dataIn[3693]),
.io_dataIn_3694(dataIn[3694]),
.io_dataIn_3695(dataIn[3695]),
.io_dataIn_3696(dataIn[3696]),
.io_dataIn_3697(dataIn[3697]),
.io_dataIn_3698(dataIn[3698]),
.io_dataIn_3699(dataIn[3699]),
.io_dataIn_3700(dataIn[3700]),
.io_dataIn_3701(dataIn[3701]),
.io_dataIn_3702(dataIn[3702]),
.io_dataIn_3703(dataIn[3703]),
.io_dataIn_3704(dataIn[3704]),
.io_dataIn_3705(dataIn[3705]),
.io_dataIn_3706(dataIn[3706]),
.io_dataIn_3707(dataIn[3707]),
.io_dataIn_3708(dataIn[3708]),
.io_dataIn_3709(dataIn[3709]),
.io_dataIn_3710(dataIn[3710]),
.io_dataIn_3711(dataIn[3711]),
.io_dataIn_3712(dataIn[3712]),
.io_dataIn_3713(dataIn[3713]),
.io_dataIn_3714(dataIn[3714]),
.io_dataIn_3715(dataIn[3715]),
.io_dataIn_3716(dataIn[3716]),
.io_dataIn_3717(dataIn[3717]),
.io_dataIn_3718(dataIn[3718]),
.io_dataIn_3719(dataIn[3719]),
.io_dataIn_3720(dataIn[3720]),
.io_dataIn_3721(dataIn[3721]),
.io_dataIn_3722(dataIn[3722]),
.io_dataIn_3723(dataIn[3723]),
.io_dataIn_3724(dataIn[3724]),
.io_dataIn_3725(dataIn[3725]),
.io_dataIn_3726(dataIn[3726]),
.io_dataIn_3727(dataIn[3727]),
.io_dataIn_3728(dataIn[3728]),
.io_dataIn_3729(dataIn[3729]),
.io_dataIn_3730(dataIn[3730]),
.io_dataIn_3731(dataIn[3731]),
.io_dataIn_3732(dataIn[3732]),
.io_dataIn_3733(dataIn[3733]),
.io_dataIn_3734(dataIn[3734]),
.io_dataIn_3735(dataIn[3735]),
.io_dataIn_3736(dataIn[3736]),
.io_dataIn_3737(dataIn[3737]),
.io_dataIn_3738(dataIn[3738]),
.io_dataIn_3739(dataIn[3739]),
.io_dataIn_3740(dataIn[3740]),
.io_dataIn_3741(dataIn[3741]),
.io_dataIn_3742(dataIn[3742]),
.io_dataIn_3743(dataIn[3743]),
.io_dataIn_3744(dataIn[3744]),
.io_dataIn_3745(dataIn[3745]),
.io_dataIn_3746(dataIn[3746]),
.io_dataIn_3747(dataIn[3747]),
.io_dataIn_3748(dataIn[3748]),
.io_dataIn_3749(dataIn[3749]),
.io_dataIn_3750(dataIn[3750]),
.io_dataIn_3751(dataIn[3751]),
.io_dataIn_3752(dataIn[3752]),
.io_dataIn_3753(dataIn[3753]),
.io_dataIn_3754(dataIn[3754]),
.io_dataIn_3755(dataIn[3755]),
.io_dataIn_3756(dataIn[3756]),
.io_dataIn_3757(dataIn[3757]),
.io_dataIn_3758(dataIn[3758]),
.io_dataIn_3759(dataIn[3759]),
.io_dataIn_3760(dataIn[3760]),
.io_dataIn_3761(dataIn[3761]),
.io_dataIn_3762(dataIn[3762]),
.io_dataIn_3763(dataIn[3763]),
.io_dataIn_3764(dataIn[3764]),
.io_dataIn_3765(dataIn[3765]),
.io_dataIn_3766(dataIn[3766]),
.io_dataIn_3767(dataIn[3767]),
.io_dataIn_3768(dataIn[3768]),
.io_dataIn_3769(dataIn[3769]),
.io_dataIn_3770(dataIn[3770]),
.io_dataIn_3771(dataIn[3771]),
.io_dataIn_3772(dataIn[3772]),
.io_dataIn_3773(dataIn[3773]),
.io_dataIn_3774(dataIn[3774]),
.io_dataIn_3775(dataIn[3775]),
.io_dataIn_3776(dataIn[3776]),
.io_dataIn_3777(dataIn[3777]),
.io_dataIn_3778(dataIn[3778]),
.io_dataIn_3779(dataIn[3779]),
.io_dataIn_3780(dataIn[3780]),
.io_dataIn_3781(dataIn[3781]),
.io_dataIn_3782(dataIn[3782]),
.io_dataIn_3783(dataIn[3783]),
.io_dataIn_3784(dataIn[3784]),
.io_dataIn_3785(dataIn[3785]),
.io_dataIn_3786(dataIn[3786]),
.io_dataIn_3787(dataIn[3787]),
.io_dataIn_3788(dataIn[3788]),
.io_dataIn_3789(dataIn[3789]),
.io_dataIn_3790(dataIn[3790]),
.io_dataIn_3791(dataIn[3791]),
.io_dataIn_3792(dataIn[3792]),
.io_dataIn_3793(dataIn[3793]),
.io_dataIn_3794(dataIn[3794]),
.io_dataIn_3795(dataIn[3795]),
.io_dataIn_3796(dataIn[3796]),
.io_dataIn_3797(dataIn[3797]),
.io_dataIn_3798(dataIn[3798]),
.io_dataIn_3799(dataIn[3799]),
.io_dataIn_3800(dataIn[3800]),
.io_dataIn_3801(dataIn[3801]),
.io_dataIn_3802(dataIn[3802]),
.io_dataIn_3803(dataIn[3803]),
.io_dataIn_3804(dataIn[3804]),
.io_dataIn_3805(dataIn[3805]),
.io_dataIn_3806(dataIn[3806]),
.io_dataIn_3807(dataIn[3807]),
.io_dataIn_3808(dataIn[3808]),
.io_dataIn_3809(dataIn[3809]),
.io_dataIn_3810(dataIn[3810]),
.io_dataIn_3811(dataIn[3811]),
.io_dataIn_3812(dataIn[3812]),
.io_dataIn_3813(dataIn[3813]),
.io_dataIn_3814(dataIn[3814]),
.io_dataIn_3815(dataIn[3815]),
.io_dataIn_3816(dataIn[3816]),
.io_dataIn_3817(dataIn[3817]),
.io_dataIn_3818(dataIn[3818]),
.io_dataIn_3819(dataIn[3819]),
.io_dataIn_3820(dataIn[3820]),
.io_dataIn_3821(dataIn[3821]),
.io_dataIn_3822(dataIn[3822]),
.io_dataIn_3823(dataIn[3823]),
.io_dataIn_3824(dataIn[3824]),
.io_dataIn_3825(dataIn[3825]),
.io_dataIn_3826(dataIn[3826]),
.io_dataIn_3827(dataIn[3827]),
.io_dataIn_3828(dataIn[3828]),
.io_dataIn_3829(dataIn[3829]),
.io_dataIn_3830(dataIn[3830]),
.io_dataIn_3831(dataIn[3831]),
.io_dataIn_3832(dataIn[3832]),
.io_dataIn_3833(dataIn[3833]),
.io_dataIn_3834(dataIn[3834]),
.io_dataIn_3835(dataIn[3835]),
.io_dataIn_3836(dataIn[3836]),
.io_dataIn_3837(dataIn[3837]),
.io_dataIn_3838(dataIn[3838]),
.io_dataIn_3839(dataIn[3839]),
.io_dataIn_3840(dataIn[3840]),
.io_dataIn_3841(dataIn[3841]),
.io_dataIn_3842(dataIn[3842]),
.io_dataIn_3843(dataIn[3843]),
.io_dataIn_3844(dataIn[3844]),
.io_dataIn_3845(dataIn[3845]),
.io_dataIn_3846(dataIn[3846]),
.io_dataIn_3847(dataIn[3847]),
.io_dataIn_3848(dataIn[3848]),
.io_dataIn_3849(dataIn[3849]),
.io_dataIn_3850(dataIn[3850]),
.io_dataIn_3851(dataIn[3851]),
.io_dataIn_3852(dataIn[3852]),
.io_dataIn_3853(dataIn[3853]),
.io_dataIn_3854(dataIn[3854]),
.io_dataIn_3855(dataIn[3855]),
.io_dataIn_3856(dataIn[3856]),
.io_dataIn_3857(dataIn[3857]),
.io_dataIn_3858(dataIn[3858]),
.io_dataIn_3859(dataIn[3859]),
.io_dataIn_3860(dataIn[3860]),
.io_dataIn_3861(dataIn[3861]),
.io_dataIn_3862(dataIn[3862]),
.io_dataIn_3863(dataIn[3863]),
.io_dataIn_3864(dataIn[3864]),
.io_dataIn_3865(dataIn[3865]),
.io_dataIn_3866(dataIn[3866]),
.io_dataIn_3867(dataIn[3867]),
.io_dataIn_3868(dataIn[3868]),
.io_dataIn_3869(dataIn[3869]),
.io_dataIn_3870(dataIn[3870]),
.io_dataIn_3871(dataIn[3871]),
.io_dataIn_3872(dataIn[3872]),
.io_dataIn_3873(dataIn[3873]),
.io_dataIn_3874(dataIn[3874]),
.io_dataIn_3875(dataIn[3875]),
.io_dataIn_3876(dataIn[3876]),
.io_dataIn_3877(dataIn[3877]),
.io_dataIn_3878(dataIn[3878]),
.io_dataIn_3879(dataIn[3879]),
.io_dataIn_3880(dataIn[3880]),
.io_dataIn_3881(dataIn[3881]),
.io_dataIn_3882(dataIn[3882]),
.io_dataIn_3883(dataIn[3883]),
.io_dataIn_3884(dataIn[3884]),
.io_dataIn_3885(dataIn[3885]),
.io_dataIn_3886(dataIn[3886]),
.io_dataIn_3887(dataIn[3887]),
.io_dataIn_3888(dataIn[3888]),
.io_dataIn_3889(dataIn[3889]),
.io_dataIn_3890(dataIn[3890]),
.io_dataIn_3891(dataIn[3891]),
.io_dataIn_3892(dataIn[3892]),
.io_dataIn_3893(dataIn[3893]),
.io_dataIn_3894(dataIn[3894]),
.io_dataIn_3895(dataIn[3895]),
.io_dataIn_3896(dataIn[3896]),
.io_dataIn_3897(dataIn[3897]),
.io_dataIn_3898(dataIn[3898]),
.io_dataIn_3899(dataIn[3899]),
.io_dataIn_3900(dataIn[3900]),
.io_dataIn_3901(dataIn[3901]),
.io_dataIn_3902(dataIn[3902]),
.io_dataIn_3903(dataIn[3903]),
.io_dataIn_3904(dataIn[3904]),
.io_dataIn_3905(dataIn[3905]),
.io_dataIn_3906(dataIn[3906]),
.io_dataIn_3907(dataIn[3907]),
.io_dataIn_3908(dataIn[3908]),
.io_dataIn_3909(dataIn[3909]),
.io_dataIn_3910(dataIn[3910]),
.io_dataIn_3911(dataIn[3911]),
.io_dataIn_3912(dataIn[3912]),
.io_dataIn_3913(dataIn[3913]),
.io_dataIn_3914(dataIn[3914]),
.io_dataIn_3915(dataIn[3915]),
.io_dataIn_3916(dataIn[3916]),
.io_dataIn_3917(dataIn[3917]),
.io_dataIn_3918(dataIn[3918]),
.io_dataIn_3919(dataIn[3919]),
.io_dataIn_3920(dataIn[3920]),
.io_dataIn_3921(dataIn[3921]),
.io_dataIn_3922(dataIn[3922]),
.io_dataIn_3923(dataIn[3923]),
.io_dataIn_3924(dataIn[3924]),
.io_dataIn_3925(dataIn[3925]),
.io_dataIn_3926(dataIn[3926]),
.io_dataIn_3927(dataIn[3927]),
.io_dataIn_3928(dataIn[3928]),
.io_dataIn_3929(dataIn[3929]),
.io_dataIn_3930(dataIn[3930]),
.io_dataIn_3931(dataIn[3931]),
.io_dataIn_3932(dataIn[3932]),
.io_dataIn_3933(dataIn[3933]),
.io_dataIn_3934(dataIn[3934]),
.io_dataIn_3935(dataIn[3935]),
.io_dataIn_3936(dataIn[3936]),
.io_dataIn_3937(dataIn[3937]),
.io_dataIn_3938(dataIn[3938]),
.io_dataIn_3939(dataIn[3939]),
.io_dataIn_3940(dataIn[3940]),
.io_dataIn_3941(dataIn[3941]),
.io_dataIn_3942(dataIn[3942]),
.io_dataIn_3943(dataIn[3943]),
.io_dataIn_3944(dataIn[3944]),
.io_dataIn_3945(dataIn[3945]),
.io_dataIn_3946(dataIn[3946]),
.io_dataIn_3947(dataIn[3947]),
.io_dataIn_3948(dataIn[3948]),
.io_dataIn_3949(dataIn[3949]),
.io_dataIn_3950(dataIn[3950]),
.io_dataIn_3951(dataIn[3951]),
.io_dataIn_3952(dataIn[3952]),
.io_dataIn_3953(dataIn[3953]),
.io_dataIn_3954(dataIn[3954]),
.io_dataIn_3955(dataIn[3955]),
.io_dataIn_3956(dataIn[3956]),
.io_dataIn_3957(dataIn[3957]),
.io_dataIn_3958(dataIn[3958]),
.io_dataIn_3959(dataIn[3959]),
.io_dataIn_3960(dataIn[3960]),
.io_dataIn_3961(dataIn[3961]),
.io_dataIn_3962(dataIn[3962]),
.io_dataIn_3963(dataIn[3963]),
.io_dataIn_3964(dataIn[3964]),
.io_dataIn_3965(dataIn[3965]),
.io_dataIn_3966(dataIn[3966]),
.io_dataIn_3967(dataIn[3967]),
.io_dataIn_3968(dataIn[3968]),
.io_dataIn_3969(dataIn[3969]),
.io_dataIn_3970(dataIn[3970]),
.io_dataIn_3971(dataIn[3971]),
.io_dataIn_3972(dataIn[3972]),
.io_dataIn_3973(dataIn[3973]),
.io_dataIn_3974(dataIn[3974]),
.io_dataIn_3975(dataIn[3975]),
.io_dataIn_3976(dataIn[3976]),
.io_dataIn_3977(dataIn[3977]),
.io_dataIn_3978(dataIn[3978]),
.io_dataIn_3979(dataIn[3979]),
.io_dataIn_3980(dataIn[3980]),
.io_dataIn_3981(dataIn[3981]),
.io_dataIn_3982(dataIn[3982]),
.io_dataIn_3983(dataIn[3983]),
.io_dataIn_3984(dataIn[3984]),
.io_dataIn_3985(dataIn[3985]),
.io_dataIn_3986(dataIn[3986]),
.io_dataIn_3987(dataIn[3987]),
.io_dataIn_3988(dataIn[3988]),
.io_dataIn_3989(dataIn[3989]),
.io_dataIn_3990(dataIn[3990]),
.io_dataIn_3991(dataIn[3991]),
.io_dataIn_3992(dataIn[3992]),
.io_dataIn_3993(dataIn[3993]),
.io_dataIn_3994(dataIn[3994]),
.io_dataIn_3995(dataIn[3995]),
.io_dataIn_3996(dataIn[3996]),
.io_dataIn_3997(dataIn[3997]),
.io_dataIn_3998(dataIn[3998]),
.io_dataIn_3999(dataIn[3999]),
.io_dataIn_4000(dataIn[4000]),
.io_dataIn_4001(dataIn[4001]),
.io_dataIn_4002(dataIn[4002]),
.io_dataIn_4003(dataIn[4003]),
.io_dataIn_4004(dataIn[4004]),
.io_dataIn_4005(dataIn[4005]),
.io_dataIn_4006(dataIn[4006]),
.io_dataIn_4007(dataIn[4007]),
.io_dataIn_4008(dataIn[4008]),
.io_dataIn_4009(dataIn[4009]),
.io_dataIn_4010(dataIn[4010]),
.io_dataIn_4011(dataIn[4011]),
.io_dataIn_4012(dataIn[4012]),
.io_dataIn_4013(dataIn[4013]),
.io_dataIn_4014(dataIn[4014]),
.io_dataIn_4015(dataIn[4015]),
.io_dataIn_4016(dataIn[4016]),
.io_dataIn_4017(dataIn[4017]),
.io_dataIn_4018(dataIn[4018]),
.io_dataIn_4019(dataIn[4019]),
.io_dataIn_4020(dataIn[4020]),
.io_dataIn_4021(dataIn[4021]),
.io_dataIn_4022(dataIn[4022]),
.io_dataIn_4023(dataIn[4023]),
.io_dataIn_4024(dataIn[4024]),
.io_dataIn_4025(dataIn[4025]),
.io_dataIn_4026(dataIn[4026]),
.io_dataIn_4027(dataIn[4027]),
.io_dataIn_4028(dataIn[4028]),
.io_dataIn_4029(dataIn[4029]),
.io_dataIn_4030(dataIn[4030]),
.io_dataIn_4031(dataIn[4031]),
.io_dataIn_4032(dataIn[4032]),
.io_dataIn_4033(dataIn[4033]),
.io_dataIn_4034(dataIn[4034]),
.io_dataIn_4035(dataIn[4035]),
.io_dataIn_4036(dataIn[4036]),
.io_dataIn_4037(dataIn[4037]),
.io_dataIn_4038(dataIn[4038]),
.io_dataIn_4039(dataIn[4039]),
.io_dataIn_4040(dataIn[4040]),
.io_dataIn_4041(dataIn[4041]),
.io_dataIn_4042(dataIn[4042]),
.io_dataIn_4043(dataIn[4043]),
.io_dataIn_4044(dataIn[4044]),
.io_dataIn_4045(dataIn[4045]),
.io_dataIn_4046(dataIn[4046]),
.io_dataIn_4047(dataIn[4047]),
.io_dataIn_4048(dataIn[4048]),
.io_dataIn_4049(dataIn[4049]),
.io_dataIn_4050(dataIn[4050]),
.io_dataIn_4051(dataIn[4051]),
.io_dataIn_4052(dataIn[4052]),
.io_dataIn_4053(dataIn[4053]),
.io_dataIn_4054(dataIn[4054]),
.io_dataIn_4055(dataIn[4055]),
.io_dataIn_4056(dataIn[4056]),
.io_dataIn_4057(dataIn[4057]),
.io_dataIn_4058(dataIn[4058]),
.io_dataIn_4059(dataIn[4059]),
.io_dataIn_4060(dataIn[4060]),
.io_dataIn_4061(dataIn[4061]),
.io_dataIn_4062(dataIn[4062]),
.io_dataIn_4063(dataIn[4063]),
.io_dataIn_4064(dataIn[4064]),
.io_dataIn_4065(dataIn[4065]),
.io_dataIn_4066(dataIn[4066]),
.io_dataIn_4067(dataIn[4067]),
.io_dataIn_4068(dataIn[4068]),
.io_dataIn_4069(dataIn[4069]),
.io_dataIn_4070(dataIn[4070]),
.io_dataIn_4071(dataIn[4071]),
.io_dataIn_4072(dataIn[4072]),
.io_dataIn_4073(dataIn[4073]),
.io_dataIn_4074(dataIn[4074]),
.io_dataIn_4075(dataIn[4075]),
.io_dataIn_4076(dataIn[4076]),
.io_dataIn_4077(dataIn[4077]),
.io_dataIn_4078(dataIn[4078]),
.io_dataIn_4079(dataIn[4079]),
.io_dataIn_4080(dataIn[4080]),
.io_dataIn_4081(dataIn[4081]),
.io_dataIn_4082(dataIn[4082]),
.io_dataIn_4083(dataIn[4083]),
.io_dataIn_4084(dataIn[4084]),
.io_dataIn_4085(dataIn[4085]),
.io_dataIn_4086(dataIn[4086]),
.io_dataIn_4087(dataIn[4087]),
.io_dataIn_4088(dataIn[4088]),
.io_dataIn_4089(dataIn[4089]),
.io_dataIn_4090(dataIn[4090]),
.io_dataIn_4091(dataIn[4091]),
.io_dataIn_4092(dataIn[4092]),
.io_dataIn_4093(dataIn[4093]),
.io_dataIn_4094(dataIn[4094]),
.io_dataIn_4095(dataIn[4095]),
.io_dataOut_0(dataOut[0]),
.io_dataOut_1(dataOut[1]),
.io_dataOut_2(dataOut[2]),
.io_dataOut_3(dataOut[3]),
.io_dataOut_4(dataOut[4]),
.io_dataOut_5(dataOut[5]),
.io_dataOut_6(dataOut[6]),
.io_dataOut_7(dataOut[7]),
.io_dataOut_8(dataOut[8]),
.io_dataOut_9(dataOut[9]),
.io_dataOut_10(dataOut[10]),
.io_dataOut_11(dataOut[11]),
.io_dataOut_12(dataOut[12]),
.io_dataOut_13(dataOut[13]),
.io_dataOut_14(dataOut[14]),
.io_dataOut_15(dataOut[15]),
.io_dataOut_16(dataOut[16]),
.io_dataOut_17(dataOut[17]),
.io_dataOut_18(dataOut[18]),
.io_dataOut_19(dataOut[19]),
.io_dataOut_20(dataOut[20]),
.io_dataOut_21(dataOut[21]),
.io_dataOut_22(dataOut[22]),
.io_dataOut_23(dataOut[23]),
.io_dataOut_24(dataOut[24]),
.io_dataOut_25(dataOut[25]),
.io_dataOut_26(dataOut[26]),
.io_dataOut_27(dataOut[27]),
.io_dataOut_28(dataOut[28]),
.io_dataOut_29(dataOut[29]),
.io_dataOut_30(dataOut[30]),
.io_dataOut_31(dataOut[31]),
.io_dataOut_32(dataOut[32]),
.io_dataOut_33(dataOut[33]),
.io_dataOut_34(dataOut[34]),
.io_dataOut_35(dataOut[35]),
.io_dataOut_36(dataOut[36]),
.io_dataOut_37(dataOut[37]),
.io_dataOut_38(dataOut[38]),
.io_dataOut_39(dataOut[39]),
.io_dataOut_40(dataOut[40]),
.io_dataOut_41(dataOut[41]),
.io_dataOut_42(dataOut[42]),
.io_dataOut_43(dataOut[43]),
.io_dataOut_44(dataOut[44]),
.io_dataOut_45(dataOut[45]),
.io_dataOut_46(dataOut[46]),
.io_dataOut_47(dataOut[47]),
.io_dataOut_48(dataOut[48]),
.io_dataOut_49(dataOut[49]),
.io_dataOut_50(dataOut[50]),
.io_dataOut_51(dataOut[51]),
.io_dataOut_52(dataOut[52]),
.io_dataOut_53(dataOut[53]),
.io_dataOut_54(dataOut[54]),
.io_dataOut_55(dataOut[55]),
.io_dataOut_56(dataOut[56]),
.io_dataOut_57(dataOut[57]),
.io_dataOut_58(dataOut[58]),
.io_dataOut_59(dataOut[59]),
.io_dataOut_60(dataOut[60]),
.io_dataOut_61(dataOut[61]),
.io_dataOut_62(dataOut[62]),
.io_dataOut_63(dataOut[63]),
.io_dataOut_64(dataOut[64]),
.io_dataOut_65(dataOut[65]),
.io_dataOut_66(dataOut[66]),
.io_dataOut_67(dataOut[67]),
.io_dataOut_68(dataOut[68]),
.io_dataOut_69(dataOut[69]),
.io_dataOut_70(dataOut[70]),
.io_dataOut_71(dataOut[71]),
.io_dataOut_72(dataOut[72]),
.io_dataOut_73(dataOut[73]),
.io_dataOut_74(dataOut[74]),
.io_dataOut_75(dataOut[75]),
.io_dataOut_76(dataOut[76]),
.io_dataOut_77(dataOut[77]),
.io_dataOut_78(dataOut[78]),
.io_dataOut_79(dataOut[79]),
.io_dataOut_80(dataOut[80]),
.io_dataOut_81(dataOut[81]),
.io_dataOut_82(dataOut[82]),
.io_dataOut_83(dataOut[83]),
.io_dataOut_84(dataOut[84]),
.io_dataOut_85(dataOut[85]),
.io_dataOut_86(dataOut[86]),
.io_dataOut_87(dataOut[87]),
.io_dataOut_88(dataOut[88]),
.io_dataOut_89(dataOut[89]),
.io_dataOut_90(dataOut[90]),
.io_dataOut_91(dataOut[91]),
.io_dataOut_92(dataOut[92]),
.io_dataOut_93(dataOut[93]),
.io_dataOut_94(dataOut[94]),
.io_dataOut_95(dataOut[95]),
.io_dataOut_96(dataOut[96]),
.io_dataOut_97(dataOut[97]),
.io_dataOut_98(dataOut[98]),
.io_dataOut_99(dataOut[99]),
.io_dataOut_100(dataOut[100]),
.io_dataOut_101(dataOut[101]),
.io_dataOut_102(dataOut[102]),
.io_dataOut_103(dataOut[103]),
.io_dataOut_104(dataOut[104]),
.io_dataOut_105(dataOut[105]),
.io_dataOut_106(dataOut[106]),
.io_dataOut_107(dataOut[107]),
.io_dataOut_108(dataOut[108]),
.io_dataOut_109(dataOut[109]),
.io_dataOut_110(dataOut[110]),
.io_dataOut_111(dataOut[111]),
.io_dataOut_112(dataOut[112]),
.io_dataOut_113(dataOut[113]),
.io_dataOut_114(dataOut[114]),
.io_dataOut_115(dataOut[115]),
.io_dataOut_116(dataOut[116]),
.io_dataOut_117(dataOut[117]),
.io_dataOut_118(dataOut[118]),
.io_dataOut_119(dataOut[119]),
.io_dataOut_120(dataOut[120]),
.io_dataOut_121(dataOut[121]),
.io_dataOut_122(dataOut[122]),
.io_dataOut_123(dataOut[123]),
.io_dataOut_124(dataOut[124]),
.io_dataOut_125(dataOut[125]),
.io_dataOut_126(dataOut[126]),
.io_dataOut_127(dataOut[127]),
.io_dataOut_128(dataOut[128]),
.io_dataOut_129(dataOut[129]),
.io_dataOut_130(dataOut[130]),
.io_dataOut_131(dataOut[131]),
.io_dataOut_132(dataOut[132]),
.io_dataOut_133(dataOut[133]),
.io_dataOut_134(dataOut[134]),
.io_dataOut_135(dataOut[135]),
.io_dataOut_136(dataOut[136]),
.io_dataOut_137(dataOut[137]),
.io_dataOut_138(dataOut[138]),
.io_dataOut_139(dataOut[139]),
.io_dataOut_140(dataOut[140]),
.io_dataOut_141(dataOut[141]),
.io_dataOut_142(dataOut[142]),
.io_dataOut_143(dataOut[143]),
.io_dataOut_144(dataOut[144]),
.io_dataOut_145(dataOut[145]),
.io_dataOut_146(dataOut[146]),
.io_dataOut_147(dataOut[147]),
.io_dataOut_148(dataOut[148]),
.io_dataOut_149(dataOut[149]),
.io_dataOut_150(dataOut[150]),
.io_dataOut_151(dataOut[151]),
.io_dataOut_152(dataOut[152]),
.io_dataOut_153(dataOut[153]),
.io_dataOut_154(dataOut[154]),
.io_dataOut_155(dataOut[155]),
.io_dataOut_156(dataOut[156]),
.io_dataOut_157(dataOut[157]),
.io_dataOut_158(dataOut[158]),
.io_dataOut_159(dataOut[159]),
.io_dataOut_160(dataOut[160]),
.io_dataOut_161(dataOut[161]),
.io_dataOut_162(dataOut[162]),
.io_dataOut_163(dataOut[163]),
.io_dataOut_164(dataOut[164]),
.io_dataOut_165(dataOut[165]),
.io_dataOut_166(dataOut[166]),
.io_dataOut_167(dataOut[167]),
.io_dataOut_168(dataOut[168]),
.io_dataOut_169(dataOut[169]),
.io_dataOut_170(dataOut[170]),
.io_dataOut_171(dataOut[171]),
.io_dataOut_172(dataOut[172]),
.io_dataOut_173(dataOut[173]),
.io_dataOut_174(dataOut[174]),
.io_dataOut_175(dataOut[175]),
.io_dataOut_176(dataOut[176]),
.io_dataOut_177(dataOut[177]),
.io_dataOut_178(dataOut[178]),
.io_dataOut_179(dataOut[179]),
.io_dataOut_180(dataOut[180]),
.io_dataOut_181(dataOut[181]),
.io_dataOut_182(dataOut[182]),
.io_dataOut_183(dataOut[183]),
.io_dataOut_184(dataOut[184]),
.io_dataOut_185(dataOut[185]),
.io_dataOut_186(dataOut[186]),
.io_dataOut_187(dataOut[187]),
.io_dataOut_188(dataOut[188]),
.io_dataOut_189(dataOut[189]),
.io_dataOut_190(dataOut[190]),
.io_dataOut_191(dataOut[191]),
.io_dataOut_192(dataOut[192]),
.io_dataOut_193(dataOut[193]),
.io_dataOut_194(dataOut[194]),
.io_dataOut_195(dataOut[195]),
.io_dataOut_196(dataOut[196]),
.io_dataOut_197(dataOut[197]),
.io_dataOut_198(dataOut[198]),
.io_dataOut_199(dataOut[199]),
.io_dataOut_200(dataOut[200]),
.io_dataOut_201(dataOut[201]),
.io_dataOut_202(dataOut[202]),
.io_dataOut_203(dataOut[203]),
.io_dataOut_204(dataOut[204]),
.io_dataOut_205(dataOut[205]),
.io_dataOut_206(dataOut[206]),
.io_dataOut_207(dataOut[207]),
.io_dataOut_208(dataOut[208]),
.io_dataOut_209(dataOut[209]),
.io_dataOut_210(dataOut[210]),
.io_dataOut_211(dataOut[211]),
.io_dataOut_212(dataOut[212]),
.io_dataOut_213(dataOut[213]),
.io_dataOut_214(dataOut[214]),
.io_dataOut_215(dataOut[215]),
.io_dataOut_216(dataOut[216]),
.io_dataOut_217(dataOut[217]),
.io_dataOut_218(dataOut[218]),
.io_dataOut_219(dataOut[219]),
.io_dataOut_220(dataOut[220]),
.io_dataOut_221(dataOut[221]),
.io_dataOut_222(dataOut[222]),
.io_dataOut_223(dataOut[223]),
.io_dataOut_224(dataOut[224]),
.io_dataOut_225(dataOut[225]),
.io_dataOut_226(dataOut[226]),
.io_dataOut_227(dataOut[227]),
.io_dataOut_228(dataOut[228]),
.io_dataOut_229(dataOut[229]),
.io_dataOut_230(dataOut[230]),
.io_dataOut_231(dataOut[231]),
.io_dataOut_232(dataOut[232]),
.io_dataOut_233(dataOut[233]),
.io_dataOut_234(dataOut[234]),
.io_dataOut_235(dataOut[235]),
.io_dataOut_236(dataOut[236]),
.io_dataOut_237(dataOut[237]),
.io_dataOut_238(dataOut[238]),
.io_dataOut_239(dataOut[239]),
.io_dataOut_240(dataOut[240]),
.io_dataOut_241(dataOut[241]),
.io_dataOut_242(dataOut[242]),
.io_dataOut_243(dataOut[243]),
.io_dataOut_244(dataOut[244]),
.io_dataOut_245(dataOut[245]),
.io_dataOut_246(dataOut[246]),
.io_dataOut_247(dataOut[247]),
.io_dataOut_248(dataOut[248]),
.io_dataOut_249(dataOut[249]),
.io_dataOut_250(dataOut[250]),
.io_dataOut_251(dataOut[251]),
.io_dataOut_252(dataOut[252]),
.io_dataOut_253(dataOut[253]),
.io_dataOut_254(dataOut[254]),
.io_dataOut_255(dataOut[255]),
.io_dataOut_256(dataOut[256]),
.io_dataOut_257(dataOut[257]),
.io_dataOut_258(dataOut[258]),
.io_dataOut_259(dataOut[259]),
.io_dataOut_260(dataOut[260]),
.io_dataOut_261(dataOut[261]),
.io_dataOut_262(dataOut[262]),
.io_dataOut_263(dataOut[263]),
.io_dataOut_264(dataOut[264]),
.io_dataOut_265(dataOut[265]),
.io_dataOut_266(dataOut[266]),
.io_dataOut_267(dataOut[267]),
.io_dataOut_268(dataOut[268]),
.io_dataOut_269(dataOut[269]),
.io_dataOut_270(dataOut[270]),
.io_dataOut_271(dataOut[271]),
.io_dataOut_272(dataOut[272]),
.io_dataOut_273(dataOut[273]),
.io_dataOut_274(dataOut[274]),
.io_dataOut_275(dataOut[275]),
.io_dataOut_276(dataOut[276]),
.io_dataOut_277(dataOut[277]),
.io_dataOut_278(dataOut[278]),
.io_dataOut_279(dataOut[279]),
.io_dataOut_280(dataOut[280]),
.io_dataOut_281(dataOut[281]),
.io_dataOut_282(dataOut[282]),
.io_dataOut_283(dataOut[283]),
.io_dataOut_284(dataOut[284]),
.io_dataOut_285(dataOut[285]),
.io_dataOut_286(dataOut[286]),
.io_dataOut_287(dataOut[287]),
.io_dataOut_288(dataOut[288]),
.io_dataOut_289(dataOut[289]),
.io_dataOut_290(dataOut[290]),
.io_dataOut_291(dataOut[291]),
.io_dataOut_292(dataOut[292]),
.io_dataOut_293(dataOut[293]),
.io_dataOut_294(dataOut[294]),
.io_dataOut_295(dataOut[295]),
.io_dataOut_296(dataOut[296]),
.io_dataOut_297(dataOut[297]),
.io_dataOut_298(dataOut[298]),
.io_dataOut_299(dataOut[299]),
.io_dataOut_300(dataOut[300]),
.io_dataOut_301(dataOut[301]),
.io_dataOut_302(dataOut[302]),
.io_dataOut_303(dataOut[303]),
.io_dataOut_304(dataOut[304]),
.io_dataOut_305(dataOut[305]),
.io_dataOut_306(dataOut[306]),
.io_dataOut_307(dataOut[307]),
.io_dataOut_308(dataOut[308]),
.io_dataOut_309(dataOut[309]),
.io_dataOut_310(dataOut[310]),
.io_dataOut_311(dataOut[311]),
.io_dataOut_312(dataOut[312]),
.io_dataOut_313(dataOut[313]),
.io_dataOut_314(dataOut[314]),
.io_dataOut_315(dataOut[315]),
.io_dataOut_316(dataOut[316]),
.io_dataOut_317(dataOut[317]),
.io_dataOut_318(dataOut[318]),
.io_dataOut_319(dataOut[319]),
.io_dataOut_320(dataOut[320]),
.io_dataOut_321(dataOut[321]),
.io_dataOut_322(dataOut[322]),
.io_dataOut_323(dataOut[323]),
.io_dataOut_324(dataOut[324]),
.io_dataOut_325(dataOut[325]),
.io_dataOut_326(dataOut[326]),
.io_dataOut_327(dataOut[327]),
.io_dataOut_328(dataOut[328]),
.io_dataOut_329(dataOut[329]),
.io_dataOut_330(dataOut[330]),
.io_dataOut_331(dataOut[331]),
.io_dataOut_332(dataOut[332]),
.io_dataOut_333(dataOut[333]),
.io_dataOut_334(dataOut[334]),
.io_dataOut_335(dataOut[335]),
.io_dataOut_336(dataOut[336]),
.io_dataOut_337(dataOut[337]),
.io_dataOut_338(dataOut[338]),
.io_dataOut_339(dataOut[339]),
.io_dataOut_340(dataOut[340]),
.io_dataOut_341(dataOut[341]),
.io_dataOut_342(dataOut[342]),
.io_dataOut_343(dataOut[343]),
.io_dataOut_344(dataOut[344]),
.io_dataOut_345(dataOut[345]),
.io_dataOut_346(dataOut[346]),
.io_dataOut_347(dataOut[347]),
.io_dataOut_348(dataOut[348]),
.io_dataOut_349(dataOut[349]),
.io_dataOut_350(dataOut[350]),
.io_dataOut_351(dataOut[351]),
.io_dataOut_352(dataOut[352]),
.io_dataOut_353(dataOut[353]),
.io_dataOut_354(dataOut[354]),
.io_dataOut_355(dataOut[355]),
.io_dataOut_356(dataOut[356]),
.io_dataOut_357(dataOut[357]),
.io_dataOut_358(dataOut[358]),
.io_dataOut_359(dataOut[359]),
.io_dataOut_360(dataOut[360]),
.io_dataOut_361(dataOut[361]),
.io_dataOut_362(dataOut[362]),
.io_dataOut_363(dataOut[363]),
.io_dataOut_364(dataOut[364]),
.io_dataOut_365(dataOut[365]),
.io_dataOut_366(dataOut[366]),
.io_dataOut_367(dataOut[367]),
.io_dataOut_368(dataOut[368]),
.io_dataOut_369(dataOut[369]),
.io_dataOut_370(dataOut[370]),
.io_dataOut_371(dataOut[371]),
.io_dataOut_372(dataOut[372]),
.io_dataOut_373(dataOut[373]),
.io_dataOut_374(dataOut[374]),
.io_dataOut_375(dataOut[375]),
.io_dataOut_376(dataOut[376]),
.io_dataOut_377(dataOut[377]),
.io_dataOut_378(dataOut[378]),
.io_dataOut_379(dataOut[379]),
.io_dataOut_380(dataOut[380]),
.io_dataOut_381(dataOut[381]),
.io_dataOut_382(dataOut[382]),
.io_dataOut_383(dataOut[383]),
.io_dataOut_384(dataOut[384]),
.io_dataOut_385(dataOut[385]),
.io_dataOut_386(dataOut[386]),
.io_dataOut_387(dataOut[387]),
.io_dataOut_388(dataOut[388]),
.io_dataOut_389(dataOut[389]),
.io_dataOut_390(dataOut[390]),
.io_dataOut_391(dataOut[391]),
.io_dataOut_392(dataOut[392]),
.io_dataOut_393(dataOut[393]),
.io_dataOut_394(dataOut[394]),
.io_dataOut_395(dataOut[395]),
.io_dataOut_396(dataOut[396]),
.io_dataOut_397(dataOut[397]),
.io_dataOut_398(dataOut[398]),
.io_dataOut_399(dataOut[399]),
.io_dataOut_400(dataOut[400]),
.io_dataOut_401(dataOut[401]),
.io_dataOut_402(dataOut[402]),
.io_dataOut_403(dataOut[403]),
.io_dataOut_404(dataOut[404]),
.io_dataOut_405(dataOut[405]),
.io_dataOut_406(dataOut[406]),
.io_dataOut_407(dataOut[407]),
.io_dataOut_408(dataOut[408]),
.io_dataOut_409(dataOut[409]),
.io_dataOut_410(dataOut[410]),
.io_dataOut_411(dataOut[411]),
.io_dataOut_412(dataOut[412]),
.io_dataOut_413(dataOut[413]),
.io_dataOut_414(dataOut[414]),
.io_dataOut_415(dataOut[415]),
.io_dataOut_416(dataOut[416]),
.io_dataOut_417(dataOut[417]),
.io_dataOut_418(dataOut[418]),
.io_dataOut_419(dataOut[419]),
.io_dataOut_420(dataOut[420]),
.io_dataOut_421(dataOut[421]),
.io_dataOut_422(dataOut[422]),
.io_dataOut_423(dataOut[423]),
.io_dataOut_424(dataOut[424]),
.io_dataOut_425(dataOut[425]),
.io_dataOut_426(dataOut[426]),
.io_dataOut_427(dataOut[427]),
.io_dataOut_428(dataOut[428]),
.io_dataOut_429(dataOut[429]),
.io_dataOut_430(dataOut[430]),
.io_dataOut_431(dataOut[431]),
.io_dataOut_432(dataOut[432]),
.io_dataOut_433(dataOut[433]),
.io_dataOut_434(dataOut[434]),
.io_dataOut_435(dataOut[435]),
.io_dataOut_436(dataOut[436]),
.io_dataOut_437(dataOut[437]),
.io_dataOut_438(dataOut[438]),
.io_dataOut_439(dataOut[439]),
.io_dataOut_440(dataOut[440]),
.io_dataOut_441(dataOut[441]),
.io_dataOut_442(dataOut[442]),
.io_dataOut_443(dataOut[443]),
.io_dataOut_444(dataOut[444]),
.io_dataOut_445(dataOut[445]),
.io_dataOut_446(dataOut[446]),
.io_dataOut_447(dataOut[447]),
.io_dataOut_448(dataOut[448]),
.io_dataOut_449(dataOut[449]),
.io_dataOut_450(dataOut[450]),
.io_dataOut_451(dataOut[451]),
.io_dataOut_452(dataOut[452]),
.io_dataOut_453(dataOut[453]),
.io_dataOut_454(dataOut[454]),
.io_dataOut_455(dataOut[455]),
.io_dataOut_456(dataOut[456]),
.io_dataOut_457(dataOut[457]),
.io_dataOut_458(dataOut[458]),
.io_dataOut_459(dataOut[459]),
.io_dataOut_460(dataOut[460]),
.io_dataOut_461(dataOut[461]),
.io_dataOut_462(dataOut[462]),
.io_dataOut_463(dataOut[463]),
.io_dataOut_464(dataOut[464]),
.io_dataOut_465(dataOut[465]),
.io_dataOut_466(dataOut[466]),
.io_dataOut_467(dataOut[467]),
.io_dataOut_468(dataOut[468]),
.io_dataOut_469(dataOut[469]),
.io_dataOut_470(dataOut[470]),
.io_dataOut_471(dataOut[471]),
.io_dataOut_472(dataOut[472]),
.io_dataOut_473(dataOut[473]),
.io_dataOut_474(dataOut[474]),
.io_dataOut_475(dataOut[475]),
.io_dataOut_476(dataOut[476]),
.io_dataOut_477(dataOut[477]),
.io_dataOut_478(dataOut[478]),
.io_dataOut_479(dataOut[479]),
.io_dataOut_480(dataOut[480]),
.io_dataOut_481(dataOut[481]),
.io_dataOut_482(dataOut[482]),
.io_dataOut_483(dataOut[483]),
.io_dataOut_484(dataOut[484]),
.io_dataOut_485(dataOut[485]),
.io_dataOut_486(dataOut[486]),
.io_dataOut_487(dataOut[487]),
.io_dataOut_488(dataOut[488]),
.io_dataOut_489(dataOut[489]),
.io_dataOut_490(dataOut[490]),
.io_dataOut_491(dataOut[491]),
.io_dataOut_492(dataOut[492]),
.io_dataOut_493(dataOut[493]),
.io_dataOut_494(dataOut[494]),
.io_dataOut_495(dataOut[495]),
.io_dataOut_496(dataOut[496]),
.io_dataOut_497(dataOut[497]),
.io_dataOut_498(dataOut[498]),
.io_dataOut_499(dataOut[499]),
.io_dataOut_500(dataOut[500]),
.io_dataOut_501(dataOut[501]),
.io_dataOut_502(dataOut[502]),
.io_dataOut_503(dataOut[503]),
.io_dataOut_504(dataOut[504]),
.io_dataOut_505(dataOut[505]),
.io_dataOut_506(dataOut[506]),
.io_dataOut_507(dataOut[507]),
.io_dataOut_508(dataOut[508]),
.io_dataOut_509(dataOut[509]),
.io_dataOut_510(dataOut[510]),
.io_dataOut_511(dataOut[511]),
.io_dataOut_512(dataOut[512]),
.io_dataOut_513(dataOut[513]),
.io_dataOut_514(dataOut[514]),
.io_dataOut_515(dataOut[515]),
.io_dataOut_516(dataOut[516]),
.io_dataOut_517(dataOut[517]),
.io_dataOut_518(dataOut[518]),
.io_dataOut_519(dataOut[519]),
.io_dataOut_520(dataOut[520]),
.io_dataOut_521(dataOut[521]),
.io_dataOut_522(dataOut[522]),
.io_dataOut_523(dataOut[523]),
.io_dataOut_524(dataOut[524]),
.io_dataOut_525(dataOut[525]),
.io_dataOut_526(dataOut[526]),
.io_dataOut_527(dataOut[527]),
.io_dataOut_528(dataOut[528]),
.io_dataOut_529(dataOut[529]),
.io_dataOut_530(dataOut[530]),
.io_dataOut_531(dataOut[531]),
.io_dataOut_532(dataOut[532]),
.io_dataOut_533(dataOut[533]),
.io_dataOut_534(dataOut[534]),
.io_dataOut_535(dataOut[535]),
.io_dataOut_536(dataOut[536]),
.io_dataOut_537(dataOut[537]),
.io_dataOut_538(dataOut[538]),
.io_dataOut_539(dataOut[539]),
.io_dataOut_540(dataOut[540]),
.io_dataOut_541(dataOut[541]),
.io_dataOut_542(dataOut[542]),
.io_dataOut_543(dataOut[543]),
.io_dataOut_544(dataOut[544]),
.io_dataOut_545(dataOut[545]),
.io_dataOut_546(dataOut[546]),
.io_dataOut_547(dataOut[547]),
.io_dataOut_548(dataOut[548]),
.io_dataOut_549(dataOut[549]),
.io_dataOut_550(dataOut[550]),
.io_dataOut_551(dataOut[551]),
.io_dataOut_552(dataOut[552]),
.io_dataOut_553(dataOut[553]),
.io_dataOut_554(dataOut[554]),
.io_dataOut_555(dataOut[555]),
.io_dataOut_556(dataOut[556]),
.io_dataOut_557(dataOut[557]),
.io_dataOut_558(dataOut[558]),
.io_dataOut_559(dataOut[559]),
.io_dataOut_560(dataOut[560]),
.io_dataOut_561(dataOut[561]),
.io_dataOut_562(dataOut[562]),
.io_dataOut_563(dataOut[563]),
.io_dataOut_564(dataOut[564]),
.io_dataOut_565(dataOut[565]),
.io_dataOut_566(dataOut[566]),
.io_dataOut_567(dataOut[567]),
.io_dataOut_568(dataOut[568]),
.io_dataOut_569(dataOut[569]),
.io_dataOut_570(dataOut[570]),
.io_dataOut_571(dataOut[571]),
.io_dataOut_572(dataOut[572]),
.io_dataOut_573(dataOut[573]),
.io_dataOut_574(dataOut[574]),
.io_dataOut_575(dataOut[575]),
.io_dataOut_576(dataOut[576]),
.io_dataOut_577(dataOut[577]),
.io_dataOut_578(dataOut[578]),
.io_dataOut_579(dataOut[579]),
.io_dataOut_580(dataOut[580]),
.io_dataOut_581(dataOut[581]),
.io_dataOut_582(dataOut[582]),
.io_dataOut_583(dataOut[583]),
.io_dataOut_584(dataOut[584]),
.io_dataOut_585(dataOut[585]),
.io_dataOut_586(dataOut[586]),
.io_dataOut_587(dataOut[587]),
.io_dataOut_588(dataOut[588]),
.io_dataOut_589(dataOut[589]),
.io_dataOut_590(dataOut[590]),
.io_dataOut_591(dataOut[591]),
.io_dataOut_592(dataOut[592]),
.io_dataOut_593(dataOut[593]),
.io_dataOut_594(dataOut[594]),
.io_dataOut_595(dataOut[595]),
.io_dataOut_596(dataOut[596]),
.io_dataOut_597(dataOut[597]),
.io_dataOut_598(dataOut[598]),
.io_dataOut_599(dataOut[599]),
.io_dataOut_600(dataOut[600]),
.io_dataOut_601(dataOut[601]),
.io_dataOut_602(dataOut[602]),
.io_dataOut_603(dataOut[603]),
.io_dataOut_604(dataOut[604]),
.io_dataOut_605(dataOut[605]),
.io_dataOut_606(dataOut[606]),
.io_dataOut_607(dataOut[607]),
.io_dataOut_608(dataOut[608]),
.io_dataOut_609(dataOut[609]),
.io_dataOut_610(dataOut[610]),
.io_dataOut_611(dataOut[611]),
.io_dataOut_612(dataOut[612]),
.io_dataOut_613(dataOut[613]),
.io_dataOut_614(dataOut[614]),
.io_dataOut_615(dataOut[615]),
.io_dataOut_616(dataOut[616]),
.io_dataOut_617(dataOut[617]),
.io_dataOut_618(dataOut[618]),
.io_dataOut_619(dataOut[619]),
.io_dataOut_620(dataOut[620]),
.io_dataOut_621(dataOut[621]),
.io_dataOut_622(dataOut[622]),
.io_dataOut_623(dataOut[623]),
.io_dataOut_624(dataOut[624]),
.io_dataOut_625(dataOut[625]),
.io_dataOut_626(dataOut[626]),
.io_dataOut_627(dataOut[627]),
.io_dataOut_628(dataOut[628]),
.io_dataOut_629(dataOut[629]),
.io_dataOut_630(dataOut[630]),
.io_dataOut_631(dataOut[631]),
.io_dataOut_632(dataOut[632]),
.io_dataOut_633(dataOut[633]),
.io_dataOut_634(dataOut[634]),
.io_dataOut_635(dataOut[635]),
.io_dataOut_636(dataOut[636]),
.io_dataOut_637(dataOut[637]),
.io_dataOut_638(dataOut[638]),
.io_dataOut_639(dataOut[639]),
.io_dataOut_640(dataOut[640]),
.io_dataOut_641(dataOut[641]),
.io_dataOut_642(dataOut[642]),
.io_dataOut_643(dataOut[643]),
.io_dataOut_644(dataOut[644]),
.io_dataOut_645(dataOut[645]),
.io_dataOut_646(dataOut[646]),
.io_dataOut_647(dataOut[647]),
.io_dataOut_648(dataOut[648]),
.io_dataOut_649(dataOut[649]),
.io_dataOut_650(dataOut[650]),
.io_dataOut_651(dataOut[651]),
.io_dataOut_652(dataOut[652]),
.io_dataOut_653(dataOut[653]),
.io_dataOut_654(dataOut[654]),
.io_dataOut_655(dataOut[655]),
.io_dataOut_656(dataOut[656]),
.io_dataOut_657(dataOut[657]),
.io_dataOut_658(dataOut[658]),
.io_dataOut_659(dataOut[659]),
.io_dataOut_660(dataOut[660]),
.io_dataOut_661(dataOut[661]),
.io_dataOut_662(dataOut[662]),
.io_dataOut_663(dataOut[663]),
.io_dataOut_664(dataOut[664]),
.io_dataOut_665(dataOut[665]),
.io_dataOut_666(dataOut[666]),
.io_dataOut_667(dataOut[667]),
.io_dataOut_668(dataOut[668]),
.io_dataOut_669(dataOut[669]),
.io_dataOut_670(dataOut[670]),
.io_dataOut_671(dataOut[671]),
.io_dataOut_672(dataOut[672]),
.io_dataOut_673(dataOut[673]),
.io_dataOut_674(dataOut[674]),
.io_dataOut_675(dataOut[675]),
.io_dataOut_676(dataOut[676]),
.io_dataOut_677(dataOut[677]),
.io_dataOut_678(dataOut[678]),
.io_dataOut_679(dataOut[679]),
.io_dataOut_680(dataOut[680]),
.io_dataOut_681(dataOut[681]),
.io_dataOut_682(dataOut[682]),
.io_dataOut_683(dataOut[683]),
.io_dataOut_684(dataOut[684]),
.io_dataOut_685(dataOut[685]),
.io_dataOut_686(dataOut[686]),
.io_dataOut_687(dataOut[687]),
.io_dataOut_688(dataOut[688]),
.io_dataOut_689(dataOut[689]),
.io_dataOut_690(dataOut[690]),
.io_dataOut_691(dataOut[691]),
.io_dataOut_692(dataOut[692]),
.io_dataOut_693(dataOut[693]),
.io_dataOut_694(dataOut[694]),
.io_dataOut_695(dataOut[695]),
.io_dataOut_696(dataOut[696]),
.io_dataOut_697(dataOut[697]),
.io_dataOut_698(dataOut[698]),
.io_dataOut_699(dataOut[699]),
.io_dataOut_700(dataOut[700]),
.io_dataOut_701(dataOut[701]),
.io_dataOut_702(dataOut[702]),
.io_dataOut_703(dataOut[703]),
.io_dataOut_704(dataOut[704]),
.io_dataOut_705(dataOut[705]),
.io_dataOut_706(dataOut[706]),
.io_dataOut_707(dataOut[707]),
.io_dataOut_708(dataOut[708]),
.io_dataOut_709(dataOut[709]),
.io_dataOut_710(dataOut[710]),
.io_dataOut_711(dataOut[711]),
.io_dataOut_712(dataOut[712]),
.io_dataOut_713(dataOut[713]),
.io_dataOut_714(dataOut[714]),
.io_dataOut_715(dataOut[715]),
.io_dataOut_716(dataOut[716]),
.io_dataOut_717(dataOut[717]),
.io_dataOut_718(dataOut[718]),
.io_dataOut_719(dataOut[719]),
.io_dataOut_720(dataOut[720]),
.io_dataOut_721(dataOut[721]),
.io_dataOut_722(dataOut[722]),
.io_dataOut_723(dataOut[723]),
.io_dataOut_724(dataOut[724]),
.io_dataOut_725(dataOut[725]),
.io_dataOut_726(dataOut[726]),
.io_dataOut_727(dataOut[727]),
.io_dataOut_728(dataOut[728]),
.io_dataOut_729(dataOut[729]),
.io_dataOut_730(dataOut[730]),
.io_dataOut_731(dataOut[731]),
.io_dataOut_732(dataOut[732]),
.io_dataOut_733(dataOut[733]),
.io_dataOut_734(dataOut[734]),
.io_dataOut_735(dataOut[735]),
.io_dataOut_736(dataOut[736]),
.io_dataOut_737(dataOut[737]),
.io_dataOut_738(dataOut[738]),
.io_dataOut_739(dataOut[739]),
.io_dataOut_740(dataOut[740]),
.io_dataOut_741(dataOut[741]),
.io_dataOut_742(dataOut[742]),
.io_dataOut_743(dataOut[743]),
.io_dataOut_744(dataOut[744]),
.io_dataOut_745(dataOut[745]),
.io_dataOut_746(dataOut[746]),
.io_dataOut_747(dataOut[747]),
.io_dataOut_748(dataOut[748]),
.io_dataOut_749(dataOut[749]),
.io_dataOut_750(dataOut[750]),
.io_dataOut_751(dataOut[751]),
.io_dataOut_752(dataOut[752]),
.io_dataOut_753(dataOut[753]),
.io_dataOut_754(dataOut[754]),
.io_dataOut_755(dataOut[755]),
.io_dataOut_756(dataOut[756]),
.io_dataOut_757(dataOut[757]),
.io_dataOut_758(dataOut[758]),
.io_dataOut_759(dataOut[759]),
.io_dataOut_760(dataOut[760]),
.io_dataOut_761(dataOut[761]),
.io_dataOut_762(dataOut[762]),
.io_dataOut_763(dataOut[763]),
.io_dataOut_764(dataOut[764]),
.io_dataOut_765(dataOut[765]),
.io_dataOut_766(dataOut[766]),
.io_dataOut_767(dataOut[767]),
.io_dataOut_768(dataOut[768]),
.io_dataOut_769(dataOut[769]),
.io_dataOut_770(dataOut[770]),
.io_dataOut_771(dataOut[771]),
.io_dataOut_772(dataOut[772]),
.io_dataOut_773(dataOut[773]),
.io_dataOut_774(dataOut[774]),
.io_dataOut_775(dataOut[775]),
.io_dataOut_776(dataOut[776]),
.io_dataOut_777(dataOut[777]),
.io_dataOut_778(dataOut[778]),
.io_dataOut_779(dataOut[779]),
.io_dataOut_780(dataOut[780]),
.io_dataOut_781(dataOut[781]),
.io_dataOut_782(dataOut[782]),
.io_dataOut_783(dataOut[783]),
.io_dataOut_784(dataOut[784]),
.io_dataOut_785(dataOut[785]),
.io_dataOut_786(dataOut[786]),
.io_dataOut_787(dataOut[787]),
.io_dataOut_788(dataOut[788]),
.io_dataOut_789(dataOut[789]),
.io_dataOut_790(dataOut[790]),
.io_dataOut_791(dataOut[791]),
.io_dataOut_792(dataOut[792]),
.io_dataOut_793(dataOut[793]),
.io_dataOut_794(dataOut[794]),
.io_dataOut_795(dataOut[795]),
.io_dataOut_796(dataOut[796]),
.io_dataOut_797(dataOut[797]),
.io_dataOut_798(dataOut[798]),
.io_dataOut_799(dataOut[799]),
.io_dataOut_800(dataOut[800]),
.io_dataOut_801(dataOut[801]),
.io_dataOut_802(dataOut[802]),
.io_dataOut_803(dataOut[803]),
.io_dataOut_804(dataOut[804]),
.io_dataOut_805(dataOut[805]),
.io_dataOut_806(dataOut[806]),
.io_dataOut_807(dataOut[807]),
.io_dataOut_808(dataOut[808]),
.io_dataOut_809(dataOut[809]),
.io_dataOut_810(dataOut[810]),
.io_dataOut_811(dataOut[811]),
.io_dataOut_812(dataOut[812]),
.io_dataOut_813(dataOut[813]),
.io_dataOut_814(dataOut[814]),
.io_dataOut_815(dataOut[815]),
.io_dataOut_816(dataOut[816]),
.io_dataOut_817(dataOut[817]),
.io_dataOut_818(dataOut[818]),
.io_dataOut_819(dataOut[819]),
.io_dataOut_820(dataOut[820]),
.io_dataOut_821(dataOut[821]),
.io_dataOut_822(dataOut[822]),
.io_dataOut_823(dataOut[823]),
.io_dataOut_824(dataOut[824]),
.io_dataOut_825(dataOut[825]),
.io_dataOut_826(dataOut[826]),
.io_dataOut_827(dataOut[827]),
.io_dataOut_828(dataOut[828]),
.io_dataOut_829(dataOut[829]),
.io_dataOut_830(dataOut[830]),
.io_dataOut_831(dataOut[831]),
.io_dataOut_832(dataOut[832]),
.io_dataOut_833(dataOut[833]),
.io_dataOut_834(dataOut[834]),
.io_dataOut_835(dataOut[835]),
.io_dataOut_836(dataOut[836]),
.io_dataOut_837(dataOut[837]),
.io_dataOut_838(dataOut[838]),
.io_dataOut_839(dataOut[839]),
.io_dataOut_840(dataOut[840]),
.io_dataOut_841(dataOut[841]),
.io_dataOut_842(dataOut[842]),
.io_dataOut_843(dataOut[843]),
.io_dataOut_844(dataOut[844]),
.io_dataOut_845(dataOut[845]),
.io_dataOut_846(dataOut[846]),
.io_dataOut_847(dataOut[847]),
.io_dataOut_848(dataOut[848]),
.io_dataOut_849(dataOut[849]),
.io_dataOut_850(dataOut[850]),
.io_dataOut_851(dataOut[851]),
.io_dataOut_852(dataOut[852]),
.io_dataOut_853(dataOut[853]),
.io_dataOut_854(dataOut[854]),
.io_dataOut_855(dataOut[855]),
.io_dataOut_856(dataOut[856]),
.io_dataOut_857(dataOut[857]),
.io_dataOut_858(dataOut[858]),
.io_dataOut_859(dataOut[859]),
.io_dataOut_860(dataOut[860]),
.io_dataOut_861(dataOut[861]),
.io_dataOut_862(dataOut[862]),
.io_dataOut_863(dataOut[863]),
.io_dataOut_864(dataOut[864]),
.io_dataOut_865(dataOut[865]),
.io_dataOut_866(dataOut[866]),
.io_dataOut_867(dataOut[867]),
.io_dataOut_868(dataOut[868]),
.io_dataOut_869(dataOut[869]),
.io_dataOut_870(dataOut[870]),
.io_dataOut_871(dataOut[871]),
.io_dataOut_872(dataOut[872]),
.io_dataOut_873(dataOut[873]),
.io_dataOut_874(dataOut[874]),
.io_dataOut_875(dataOut[875]),
.io_dataOut_876(dataOut[876]),
.io_dataOut_877(dataOut[877]),
.io_dataOut_878(dataOut[878]),
.io_dataOut_879(dataOut[879]),
.io_dataOut_880(dataOut[880]),
.io_dataOut_881(dataOut[881]),
.io_dataOut_882(dataOut[882]),
.io_dataOut_883(dataOut[883]),
.io_dataOut_884(dataOut[884]),
.io_dataOut_885(dataOut[885]),
.io_dataOut_886(dataOut[886]),
.io_dataOut_887(dataOut[887]),
.io_dataOut_888(dataOut[888]),
.io_dataOut_889(dataOut[889]),
.io_dataOut_890(dataOut[890]),
.io_dataOut_891(dataOut[891]),
.io_dataOut_892(dataOut[892]),
.io_dataOut_893(dataOut[893]),
.io_dataOut_894(dataOut[894]),
.io_dataOut_895(dataOut[895]),
.io_dataOut_896(dataOut[896]),
.io_dataOut_897(dataOut[897]),
.io_dataOut_898(dataOut[898]),
.io_dataOut_899(dataOut[899]),
.io_dataOut_900(dataOut[900]),
.io_dataOut_901(dataOut[901]),
.io_dataOut_902(dataOut[902]),
.io_dataOut_903(dataOut[903]),
.io_dataOut_904(dataOut[904]),
.io_dataOut_905(dataOut[905]),
.io_dataOut_906(dataOut[906]),
.io_dataOut_907(dataOut[907]),
.io_dataOut_908(dataOut[908]),
.io_dataOut_909(dataOut[909]),
.io_dataOut_910(dataOut[910]),
.io_dataOut_911(dataOut[911]),
.io_dataOut_912(dataOut[912]),
.io_dataOut_913(dataOut[913]),
.io_dataOut_914(dataOut[914]),
.io_dataOut_915(dataOut[915]),
.io_dataOut_916(dataOut[916]),
.io_dataOut_917(dataOut[917]),
.io_dataOut_918(dataOut[918]),
.io_dataOut_919(dataOut[919]),
.io_dataOut_920(dataOut[920]),
.io_dataOut_921(dataOut[921]),
.io_dataOut_922(dataOut[922]),
.io_dataOut_923(dataOut[923]),
.io_dataOut_924(dataOut[924]),
.io_dataOut_925(dataOut[925]),
.io_dataOut_926(dataOut[926]),
.io_dataOut_927(dataOut[927]),
.io_dataOut_928(dataOut[928]),
.io_dataOut_929(dataOut[929]),
.io_dataOut_930(dataOut[930]),
.io_dataOut_931(dataOut[931]),
.io_dataOut_932(dataOut[932]),
.io_dataOut_933(dataOut[933]),
.io_dataOut_934(dataOut[934]),
.io_dataOut_935(dataOut[935]),
.io_dataOut_936(dataOut[936]),
.io_dataOut_937(dataOut[937]),
.io_dataOut_938(dataOut[938]),
.io_dataOut_939(dataOut[939]),
.io_dataOut_940(dataOut[940]),
.io_dataOut_941(dataOut[941]),
.io_dataOut_942(dataOut[942]),
.io_dataOut_943(dataOut[943]),
.io_dataOut_944(dataOut[944]),
.io_dataOut_945(dataOut[945]),
.io_dataOut_946(dataOut[946]),
.io_dataOut_947(dataOut[947]),
.io_dataOut_948(dataOut[948]),
.io_dataOut_949(dataOut[949]),
.io_dataOut_950(dataOut[950]),
.io_dataOut_951(dataOut[951]),
.io_dataOut_952(dataOut[952]),
.io_dataOut_953(dataOut[953]),
.io_dataOut_954(dataOut[954]),
.io_dataOut_955(dataOut[955]),
.io_dataOut_956(dataOut[956]),
.io_dataOut_957(dataOut[957]),
.io_dataOut_958(dataOut[958]),
.io_dataOut_959(dataOut[959]),
.io_dataOut_960(dataOut[960]),
.io_dataOut_961(dataOut[961]),
.io_dataOut_962(dataOut[962]),
.io_dataOut_963(dataOut[963]),
.io_dataOut_964(dataOut[964]),
.io_dataOut_965(dataOut[965]),
.io_dataOut_966(dataOut[966]),
.io_dataOut_967(dataOut[967]),
.io_dataOut_968(dataOut[968]),
.io_dataOut_969(dataOut[969]),
.io_dataOut_970(dataOut[970]),
.io_dataOut_971(dataOut[971]),
.io_dataOut_972(dataOut[972]),
.io_dataOut_973(dataOut[973]),
.io_dataOut_974(dataOut[974]),
.io_dataOut_975(dataOut[975]),
.io_dataOut_976(dataOut[976]),
.io_dataOut_977(dataOut[977]),
.io_dataOut_978(dataOut[978]),
.io_dataOut_979(dataOut[979]),
.io_dataOut_980(dataOut[980]),
.io_dataOut_981(dataOut[981]),
.io_dataOut_982(dataOut[982]),
.io_dataOut_983(dataOut[983]),
.io_dataOut_984(dataOut[984]),
.io_dataOut_985(dataOut[985]),
.io_dataOut_986(dataOut[986]),
.io_dataOut_987(dataOut[987]),
.io_dataOut_988(dataOut[988]),
.io_dataOut_989(dataOut[989]),
.io_dataOut_990(dataOut[990]),
.io_dataOut_991(dataOut[991]),
.io_dataOut_992(dataOut[992]),
.io_dataOut_993(dataOut[993]),
.io_dataOut_994(dataOut[994]),
.io_dataOut_995(dataOut[995]),
.io_dataOut_996(dataOut[996]),
.io_dataOut_997(dataOut[997]),
.io_dataOut_998(dataOut[998]),
.io_dataOut_999(dataOut[999]),
.io_dataOut_1000(dataOut[1000]),
.io_dataOut_1001(dataOut[1001]),
.io_dataOut_1002(dataOut[1002]),
.io_dataOut_1003(dataOut[1003]),
.io_dataOut_1004(dataOut[1004]),
.io_dataOut_1005(dataOut[1005]),
.io_dataOut_1006(dataOut[1006]),
.io_dataOut_1007(dataOut[1007]),
.io_dataOut_1008(dataOut[1008]),
.io_dataOut_1009(dataOut[1009]),
.io_dataOut_1010(dataOut[1010]),
.io_dataOut_1011(dataOut[1011]),
.io_dataOut_1012(dataOut[1012]),
.io_dataOut_1013(dataOut[1013]),
.io_dataOut_1014(dataOut[1014]),
.io_dataOut_1015(dataOut[1015]),
.io_dataOut_1016(dataOut[1016]),
.io_dataOut_1017(dataOut[1017]),
.io_dataOut_1018(dataOut[1018]),
.io_dataOut_1019(dataOut[1019]),
.io_dataOut_1020(dataOut[1020]),
.io_dataOut_1021(dataOut[1021]),
.io_dataOut_1022(dataOut[1022]),
.io_dataOut_1023(dataOut[1023]),
.io_dataOut_1024(dataOut[1024]),
.io_dataOut_1025(dataOut[1025]),
.io_dataOut_1026(dataOut[1026]),
.io_dataOut_1027(dataOut[1027]),
.io_dataOut_1028(dataOut[1028]),
.io_dataOut_1029(dataOut[1029]),
.io_dataOut_1030(dataOut[1030]),
.io_dataOut_1031(dataOut[1031]),
.io_dataOut_1032(dataOut[1032]),
.io_dataOut_1033(dataOut[1033]),
.io_dataOut_1034(dataOut[1034]),
.io_dataOut_1035(dataOut[1035]),
.io_dataOut_1036(dataOut[1036]),
.io_dataOut_1037(dataOut[1037]),
.io_dataOut_1038(dataOut[1038]),
.io_dataOut_1039(dataOut[1039]),
.io_dataOut_1040(dataOut[1040]),
.io_dataOut_1041(dataOut[1041]),
.io_dataOut_1042(dataOut[1042]),
.io_dataOut_1043(dataOut[1043]),
.io_dataOut_1044(dataOut[1044]),
.io_dataOut_1045(dataOut[1045]),
.io_dataOut_1046(dataOut[1046]),
.io_dataOut_1047(dataOut[1047]),
.io_dataOut_1048(dataOut[1048]),
.io_dataOut_1049(dataOut[1049]),
.io_dataOut_1050(dataOut[1050]),
.io_dataOut_1051(dataOut[1051]),
.io_dataOut_1052(dataOut[1052]),
.io_dataOut_1053(dataOut[1053]),
.io_dataOut_1054(dataOut[1054]),
.io_dataOut_1055(dataOut[1055]),
.io_dataOut_1056(dataOut[1056]),
.io_dataOut_1057(dataOut[1057]),
.io_dataOut_1058(dataOut[1058]),
.io_dataOut_1059(dataOut[1059]),
.io_dataOut_1060(dataOut[1060]),
.io_dataOut_1061(dataOut[1061]),
.io_dataOut_1062(dataOut[1062]),
.io_dataOut_1063(dataOut[1063]),
.io_dataOut_1064(dataOut[1064]),
.io_dataOut_1065(dataOut[1065]),
.io_dataOut_1066(dataOut[1066]),
.io_dataOut_1067(dataOut[1067]),
.io_dataOut_1068(dataOut[1068]),
.io_dataOut_1069(dataOut[1069]),
.io_dataOut_1070(dataOut[1070]),
.io_dataOut_1071(dataOut[1071]),
.io_dataOut_1072(dataOut[1072]),
.io_dataOut_1073(dataOut[1073]),
.io_dataOut_1074(dataOut[1074]),
.io_dataOut_1075(dataOut[1075]),
.io_dataOut_1076(dataOut[1076]),
.io_dataOut_1077(dataOut[1077]),
.io_dataOut_1078(dataOut[1078]),
.io_dataOut_1079(dataOut[1079]),
.io_dataOut_1080(dataOut[1080]),
.io_dataOut_1081(dataOut[1081]),
.io_dataOut_1082(dataOut[1082]),
.io_dataOut_1083(dataOut[1083]),
.io_dataOut_1084(dataOut[1084]),
.io_dataOut_1085(dataOut[1085]),
.io_dataOut_1086(dataOut[1086]),
.io_dataOut_1087(dataOut[1087]),
.io_dataOut_1088(dataOut[1088]),
.io_dataOut_1089(dataOut[1089]),
.io_dataOut_1090(dataOut[1090]),
.io_dataOut_1091(dataOut[1091]),
.io_dataOut_1092(dataOut[1092]),
.io_dataOut_1093(dataOut[1093]),
.io_dataOut_1094(dataOut[1094]),
.io_dataOut_1095(dataOut[1095]),
.io_dataOut_1096(dataOut[1096]),
.io_dataOut_1097(dataOut[1097]),
.io_dataOut_1098(dataOut[1098]),
.io_dataOut_1099(dataOut[1099]),
.io_dataOut_1100(dataOut[1100]),
.io_dataOut_1101(dataOut[1101]),
.io_dataOut_1102(dataOut[1102]),
.io_dataOut_1103(dataOut[1103]),
.io_dataOut_1104(dataOut[1104]),
.io_dataOut_1105(dataOut[1105]),
.io_dataOut_1106(dataOut[1106]),
.io_dataOut_1107(dataOut[1107]),
.io_dataOut_1108(dataOut[1108]),
.io_dataOut_1109(dataOut[1109]),
.io_dataOut_1110(dataOut[1110]),
.io_dataOut_1111(dataOut[1111]),
.io_dataOut_1112(dataOut[1112]),
.io_dataOut_1113(dataOut[1113]),
.io_dataOut_1114(dataOut[1114]),
.io_dataOut_1115(dataOut[1115]),
.io_dataOut_1116(dataOut[1116]),
.io_dataOut_1117(dataOut[1117]),
.io_dataOut_1118(dataOut[1118]),
.io_dataOut_1119(dataOut[1119]),
.io_dataOut_1120(dataOut[1120]),
.io_dataOut_1121(dataOut[1121]),
.io_dataOut_1122(dataOut[1122]),
.io_dataOut_1123(dataOut[1123]),
.io_dataOut_1124(dataOut[1124]),
.io_dataOut_1125(dataOut[1125]),
.io_dataOut_1126(dataOut[1126]),
.io_dataOut_1127(dataOut[1127]),
.io_dataOut_1128(dataOut[1128]),
.io_dataOut_1129(dataOut[1129]),
.io_dataOut_1130(dataOut[1130]),
.io_dataOut_1131(dataOut[1131]),
.io_dataOut_1132(dataOut[1132]),
.io_dataOut_1133(dataOut[1133]),
.io_dataOut_1134(dataOut[1134]),
.io_dataOut_1135(dataOut[1135]),
.io_dataOut_1136(dataOut[1136]),
.io_dataOut_1137(dataOut[1137]),
.io_dataOut_1138(dataOut[1138]),
.io_dataOut_1139(dataOut[1139]),
.io_dataOut_1140(dataOut[1140]),
.io_dataOut_1141(dataOut[1141]),
.io_dataOut_1142(dataOut[1142]),
.io_dataOut_1143(dataOut[1143]),
.io_dataOut_1144(dataOut[1144]),
.io_dataOut_1145(dataOut[1145]),
.io_dataOut_1146(dataOut[1146]),
.io_dataOut_1147(dataOut[1147]),
.io_dataOut_1148(dataOut[1148]),
.io_dataOut_1149(dataOut[1149]),
.io_dataOut_1150(dataOut[1150]),
.io_dataOut_1151(dataOut[1151]),
.io_dataOut_1152(dataOut[1152]),
.io_dataOut_1153(dataOut[1153]),
.io_dataOut_1154(dataOut[1154]),
.io_dataOut_1155(dataOut[1155]),
.io_dataOut_1156(dataOut[1156]),
.io_dataOut_1157(dataOut[1157]),
.io_dataOut_1158(dataOut[1158]),
.io_dataOut_1159(dataOut[1159]),
.io_dataOut_1160(dataOut[1160]),
.io_dataOut_1161(dataOut[1161]),
.io_dataOut_1162(dataOut[1162]),
.io_dataOut_1163(dataOut[1163]),
.io_dataOut_1164(dataOut[1164]),
.io_dataOut_1165(dataOut[1165]),
.io_dataOut_1166(dataOut[1166]),
.io_dataOut_1167(dataOut[1167]),
.io_dataOut_1168(dataOut[1168]),
.io_dataOut_1169(dataOut[1169]),
.io_dataOut_1170(dataOut[1170]),
.io_dataOut_1171(dataOut[1171]),
.io_dataOut_1172(dataOut[1172]),
.io_dataOut_1173(dataOut[1173]),
.io_dataOut_1174(dataOut[1174]),
.io_dataOut_1175(dataOut[1175]),
.io_dataOut_1176(dataOut[1176]),
.io_dataOut_1177(dataOut[1177]),
.io_dataOut_1178(dataOut[1178]),
.io_dataOut_1179(dataOut[1179]),
.io_dataOut_1180(dataOut[1180]),
.io_dataOut_1181(dataOut[1181]),
.io_dataOut_1182(dataOut[1182]),
.io_dataOut_1183(dataOut[1183]),
.io_dataOut_1184(dataOut[1184]),
.io_dataOut_1185(dataOut[1185]),
.io_dataOut_1186(dataOut[1186]),
.io_dataOut_1187(dataOut[1187]),
.io_dataOut_1188(dataOut[1188]),
.io_dataOut_1189(dataOut[1189]),
.io_dataOut_1190(dataOut[1190]),
.io_dataOut_1191(dataOut[1191]),
.io_dataOut_1192(dataOut[1192]),
.io_dataOut_1193(dataOut[1193]),
.io_dataOut_1194(dataOut[1194]),
.io_dataOut_1195(dataOut[1195]),
.io_dataOut_1196(dataOut[1196]),
.io_dataOut_1197(dataOut[1197]),
.io_dataOut_1198(dataOut[1198]),
.io_dataOut_1199(dataOut[1199]),
.io_dataOut_1200(dataOut[1200]),
.io_dataOut_1201(dataOut[1201]),
.io_dataOut_1202(dataOut[1202]),
.io_dataOut_1203(dataOut[1203]),
.io_dataOut_1204(dataOut[1204]),
.io_dataOut_1205(dataOut[1205]),
.io_dataOut_1206(dataOut[1206]),
.io_dataOut_1207(dataOut[1207]),
.io_dataOut_1208(dataOut[1208]),
.io_dataOut_1209(dataOut[1209]),
.io_dataOut_1210(dataOut[1210]),
.io_dataOut_1211(dataOut[1211]),
.io_dataOut_1212(dataOut[1212]),
.io_dataOut_1213(dataOut[1213]),
.io_dataOut_1214(dataOut[1214]),
.io_dataOut_1215(dataOut[1215]),
.io_dataOut_1216(dataOut[1216]),
.io_dataOut_1217(dataOut[1217]),
.io_dataOut_1218(dataOut[1218]),
.io_dataOut_1219(dataOut[1219]),
.io_dataOut_1220(dataOut[1220]),
.io_dataOut_1221(dataOut[1221]),
.io_dataOut_1222(dataOut[1222]),
.io_dataOut_1223(dataOut[1223]),
.io_dataOut_1224(dataOut[1224]),
.io_dataOut_1225(dataOut[1225]),
.io_dataOut_1226(dataOut[1226]),
.io_dataOut_1227(dataOut[1227]),
.io_dataOut_1228(dataOut[1228]),
.io_dataOut_1229(dataOut[1229]),
.io_dataOut_1230(dataOut[1230]),
.io_dataOut_1231(dataOut[1231]),
.io_dataOut_1232(dataOut[1232]),
.io_dataOut_1233(dataOut[1233]),
.io_dataOut_1234(dataOut[1234]),
.io_dataOut_1235(dataOut[1235]),
.io_dataOut_1236(dataOut[1236]),
.io_dataOut_1237(dataOut[1237]),
.io_dataOut_1238(dataOut[1238]),
.io_dataOut_1239(dataOut[1239]),
.io_dataOut_1240(dataOut[1240]),
.io_dataOut_1241(dataOut[1241]),
.io_dataOut_1242(dataOut[1242]),
.io_dataOut_1243(dataOut[1243]),
.io_dataOut_1244(dataOut[1244]),
.io_dataOut_1245(dataOut[1245]),
.io_dataOut_1246(dataOut[1246]),
.io_dataOut_1247(dataOut[1247]),
.io_dataOut_1248(dataOut[1248]),
.io_dataOut_1249(dataOut[1249]),
.io_dataOut_1250(dataOut[1250]),
.io_dataOut_1251(dataOut[1251]),
.io_dataOut_1252(dataOut[1252]),
.io_dataOut_1253(dataOut[1253]),
.io_dataOut_1254(dataOut[1254]),
.io_dataOut_1255(dataOut[1255]),
.io_dataOut_1256(dataOut[1256]),
.io_dataOut_1257(dataOut[1257]),
.io_dataOut_1258(dataOut[1258]),
.io_dataOut_1259(dataOut[1259]),
.io_dataOut_1260(dataOut[1260]),
.io_dataOut_1261(dataOut[1261]),
.io_dataOut_1262(dataOut[1262]),
.io_dataOut_1263(dataOut[1263]),
.io_dataOut_1264(dataOut[1264]),
.io_dataOut_1265(dataOut[1265]),
.io_dataOut_1266(dataOut[1266]),
.io_dataOut_1267(dataOut[1267]),
.io_dataOut_1268(dataOut[1268]),
.io_dataOut_1269(dataOut[1269]),
.io_dataOut_1270(dataOut[1270]),
.io_dataOut_1271(dataOut[1271]),
.io_dataOut_1272(dataOut[1272]),
.io_dataOut_1273(dataOut[1273]),
.io_dataOut_1274(dataOut[1274]),
.io_dataOut_1275(dataOut[1275]),
.io_dataOut_1276(dataOut[1276]),
.io_dataOut_1277(dataOut[1277]),
.io_dataOut_1278(dataOut[1278]),
.io_dataOut_1279(dataOut[1279]),
.io_dataOut_1280(dataOut[1280]),
.io_dataOut_1281(dataOut[1281]),
.io_dataOut_1282(dataOut[1282]),
.io_dataOut_1283(dataOut[1283]),
.io_dataOut_1284(dataOut[1284]),
.io_dataOut_1285(dataOut[1285]),
.io_dataOut_1286(dataOut[1286]),
.io_dataOut_1287(dataOut[1287]),
.io_dataOut_1288(dataOut[1288]),
.io_dataOut_1289(dataOut[1289]),
.io_dataOut_1290(dataOut[1290]),
.io_dataOut_1291(dataOut[1291]),
.io_dataOut_1292(dataOut[1292]),
.io_dataOut_1293(dataOut[1293]),
.io_dataOut_1294(dataOut[1294]),
.io_dataOut_1295(dataOut[1295]),
.io_dataOut_1296(dataOut[1296]),
.io_dataOut_1297(dataOut[1297]),
.io_dataOut_1298(dataOut[1298]),
.io_dataOut_1299(dataOut[1299]),
.io_dataOut_1300(dataOut[1300]),
.io_dataOut_1301(dataOut[1301]),
.io_dataOut_1302(dataOut[1302]),
.io_dataOut_1303(dataOut[1303]),
.io_dataOut_1304(dataOut[1304]),
.io_dataOut_1305(dataOut[1305]),
.io_dataOut_1306(dataOut[1306]),
.io_dataOut_1307(dataOut[1307]),
.io_dataOut_1308(dataOut[1308]),
.io_dataOut_1309(dataOut[1309]),
.io_dataOut_1310(dataOut[1310]),
.io_dataOut_1311(dataOut[1311]),
.io_dataOut_1312(dataOut[1312]),
.io_dataOut_1313(dataOut[1313]),
.io_dataOut_1314(dataOut[1314]),
.io_dataOut_1315(dataOut[1315]),
.io_dataOut_1316(dataOut[1316]),
.io_dataOut_1317(dataOut[1317]),
.io_dataOut_1318(dataOut[1318]),
.io_dataOut_1319(dataOut[1319]),
.io_dataOut_1320(dataOut[1320]),
.io_dataOut_1321(dataOut[1321]),
.io_dataOut_1322(dataOut[1322]),
.io_dataOut_1323(dataOut[1323]),
.io_dataOut_1324(dataOut[1324]),
.io_dataOut_1325(dataOut[1325]),
.io_dataOut_1326(dataOut[1326]),
.io_dataOut_1327(dataOut[1327]),
.io_dataOut_1328(dataOut[1328]),
.io_dataOut_1329(dataOut[1329]),
.io_dataOut_1330(dataOut[1330]),
.io_dataOut_1331(dataOut[1331]),
.io_dataOut_1332(dataOut[1332]),
.io_dataOut_1333(dataOut[1333]),
.io_dataOut_1334(dataOut[1334]),
.io_dataOut_1335(dataOut[1335]),
.io_dataOut_1336(dataOut[1336]),
.io_dataOut_1337(dataOut[1337]),
.io_dataOut_1338(dataOut[1338]),
.io_dataOut_1339(dataOut[1339]),
.io_dataOut_1340(dataOut[1340]),
.io_dataOut_1341(dataOut[1341]),
.io_dataOut_1342(dataOut[1342]),
.io_dataOut_1343(dataOut[1343]),
.io_dataOut_1344(dataOut[1344]),
.io_dataOut_1345(dataOut[1345]),
.io_dataOut_1346(dataOut[1346]),
.io_dataOut_1347(dataOut[1347]),
.io_dataOut_1348(dataOut[1348]),
.io_dataOut_1349(dataOut[1349]),
.io_dataOut_1350(dataOut[1350]),
.io_dataOut_1351(dataOut[1351]),
.io_dataOut_1352(dataOut[1352]),
.io_dataOut_1353(dataOut[1353]),
.io_dataOut_1354(dataOut[1354]),
.io_dataOut_1355(dataOut[1355]),
.io_dataOut_1356(dataOut[1356]),
.io_dataOut_1357(dataOut[1357]),
.io_dataOut_1358(dataOut[1358]),
.io_dataOut_1359(dataOut[1359]),
.io_dataOut_1360(dataOut[1360]),
.io_dataOut_1361(dataOut[1361]),
.io_dataOut_1362(dataOut[1362]),
.io_dataOut_1363(dataOut[1363]),
.io_dataOut_1364(dataOut[1364]),
.io_dataOut_1365(dataOut[1365]),
.io_dataOut_1366(dataOut[1366]),
.io_dataOut_1367(dataOut[1367]),
.io_dataOut_1368(dataOut[1368]),
.io_dataOut_1369(dataOut[1369]),
.io_dataOut_1370(dataOut[1370]),
.io_dataOut_1371(dataOut[1371]),
.io_dataOut_1372(dataOut[1372]),
.io_dataOut_1373(dataOut[1373]),
.io_dataOut_1374(dataOut[1374]),
.io_dataOut_1375(dataOut[1375]),
.io_dataOut_1376(dataOut[1376]),
.io_dataOut_1377(dataOut[1377]),
.io_dataOut_1378(dataOut[1378]),
.io_dataOut_1379(dataOut[1379]),
.io_dataOut_1380(dataOut[1380]),
.io_dataOut_1381(dataOut[1381]),
.io_dataOut_1382(dataOut[1382]),
.io_dataOut_1383(dataOut[1383]),
.io_dataOut_1384(dataOut[1384]),
.io_dataOut_1385(dataOut[1385]),
.io_dataOut_1386(dataOut[1386]),
.io_dataOut_1387(dataOut[1387]),
.io_dataOut_1388(dataOut[1388]),
.io_dataOut_1389(dataOut[1389]),
.io_dataOut_1390(dataOut[1390]),
.io_dataOut_1391(dataOut[1391]),
.io_dataOut_1392(dataOut[1392]),
.io_dataOut_1393(dataOut[1393]),
.io_dataOut_1394(dataOut[1394]),
.io_dataOut_1395(dataOut[1395]),
.io_dataOut_1396(dataOut[1396]),
.io_dataOut_1397(dataOut[1397]),
.io_dataOut_1398(dataOut[1398]),
.io_dataOut_1399(dataOut[1399]),
.io_dataOut_1400(dataOut[1400]),
.io_dataOut_1401(dataOut[1401]),
.io_dataOut_1402(dataOut[1402]),
.io_dataOut_1403(dataOut[1403]),
.io_dataOut_1404(dataOut[1404]),
.io_dataOut_1405(dataOut[1405]),
.io_dataOut_1406(dataOut[1406]),
.io_dataOut_1407(dataOut[1407]),
.io_dataOut_1408(dataOut[1408]),
.io_dataOut_1409(dataOut[1409]),
.io_dataOut_1410(dataOut[1410]),
.io_dataOut_1411(dataOut[1411]),
.io_dataOut_1412(dataOut[1412]),
.io_dataOut_1413(dataOut[1413]),
.io_dataOut_1414(dataOut[1414]),
.io_dataOut_1415(dataOut[1415]),
.io_dataOut_1416(dataOut[1416]),
.io_dataOut_1417(dataOut[1417]),
.io_dataOut_1418(dataOut[1418]),
.io_dataOut_1419(dataOut[1419]),
.io_dataOut_1420(dataOut[1420]),
.io_dataOut_1421(dataOut[1421]),
.io_dataOut_1422(dataOut[1422]),
.io_dataOut_1423(dataOut[1423]),
.io_dataOut_1424(dataOut[1424]),
.io_dataOut_1425(dataOut[1425]),
.io_dataOut_1426(dataOut[1426]),
.io_dataOut_1427(dataOut[1427]),
.io_dataOut_1428(dataOut[1428]),
.io_dataOut_1429(dataOut[1429]),
.io_dataOut_1430(dataOut[1430]),
.io_dataOut_1431(dataOut[1431]),
.io_dataOut_1432(dataOut[1432]),
.io_dataOut_1433(dataOut[1433]),
.io_dataOut_1434(dataOut[1434]),
.io_dataOut_1435(dataOut[1435]),
.io_dataOut_1436(dataOut[1436]),
.io_dataOut_1437(dataOut[1437]),
.io_dataOut_1438(dataOut[1438]),
.io_dataOut_1439(dataOut[1439]),
.io_dataOut_1440(dataOut[1440]),
.io_dataOut_1441(dataOut[1441]),
.io_dataOut_1442(dataOut[1442]),
.io_dataOut_1443(dataOut[1443]),
.io_dataOut_1444(dataOut[1444]),
.io_dataOut_1445(dataOut[1445]),
.io_dataOut_1446(dataOut[1446]),
.io_dataOut_1447(dataOut[1447]),
.io_dataOut_1448(dataOut[1448]),
.io_dataOut_1449(dataOut[1449]),
.io_dataOut_1450(dataOut[1450]),
.io_dataOut_1451(dataOut[1451]),
.io_dataOut_1452(dataOut[1452]),
.io_dataOut_1453(dataOut[1453]),
.io_dataOut_1454(dataOut[1454]),
.io_dataOut_1455(dataOut[1455]),
.io_dataOut_1456(dataOut[1456]),
.io_dataOut_1457(dataOut[1457]),
.io_dataOut_1458(dataOut[1458]),
.io_dataOut_1459(dataOut[1459]),
.io_dataOut_1460(dataOut[1460]),
.io_dataOut_1461(dataOut[1461]),
.io_dataOut_1462(dataOut[1462]),
.io_dataOut_1463(dataOut[1463]),
.io_dataOut_1464(dataOut[1464]),
.io_dataOut_1465(dataOut[1465]),
.io_dataOut_1466(dataOut[1466]),
.io_dataOut_1467(dataOut[1467]),
.io_dataOut_1468(dataOut[1468]),
.io_dataOut_1469(dataOut[1469]),
.io_dataOut_1470(dataOut[1470]),
.io_dataOut_1471(dataOut[1471]),
.io_dataOut_1472(dataOut[1472]),
.io_dataOut_1473(dataOut[1473]),
.io_dataOut_1474(dataOut[1474]),
.io_dataOut_1475(dataOut[1475]),
.io_dataOut_1476(dataOut[1476]),
.io_dataOut_1477(dataOut[1477]),
.io_dataOut_1478(dataOut[1478]),
.io_dataOut_1479(dataOut[1479]),
.io_dataOut_1480(dataOut[1480]),
.io_dataOut_1481(dataOut[1481]),
.io_dataOut_1482(dataOut[1482]),
.io_dataOut_1483(dataOut[1483]),
.io_dataOut_1484(dataOut[1484]),
.io_dataOut_1485(dataOut[1485]),
.io_dataOut_1486(dataOut[1486]),
.io_dataOut_1487(dataOut[1487]),
.io_dataOut_1488(dataOut[1488]),
.io_dataOut_1489(dataOut[1489]),
.io_dataOut_1490(dataOut[1490]),
.io_dataOut_1491(dataOut[1491]),
.io_dataOut_1492(dataOut[1492]),
.io_dataOut_1493(dataOut[1493]),
.io_dataOut_1494(dataOut[1494]),
.io_dataOut_1495(dataOut[1495]),
.io_dataOut_1496(dataOut[1496]),
.io_dataOut_1497(dataOut[1497]),
.io_dataOut_1498(dataOut[1498]),
.io_dataOut_1499(dataOut[1499]),
.io_dataOut_1500(dataOut[1500]),
.io_dataOut_1501(dataOut[1501]),
.io_dataOut_1502(dataOut[1502]),
.io_dataOut_1503(dataOut[1503]),
.io_dataOut_1504(dataOut[1504]),
.io_dataOut_1505(dataOut[1505]),
.io_dataOut_1506(dataOut[1506]),
.io_dataOut_1507(dataOut[1507]),
.io_dataOut_1508(dataOut[1508]),
.io_dataOut_1509(dataOut[1509]),
.io_dataOut_1510(dataOut[1510]),
.io_dataOut_1511(dataOut[1511]),
.io_dataOut_1512(dataOut[1512]),
.io_dataOut_1513(dataOut[1513]),
.io_dataOut_1514(dataOut[1514]),
.io_dataOut_1515(dataOut[1515]),
.io_dataOut_1516(dataOut[1516]),
.io_dataOut_1517(dataOut[1517]),
.io_dataOut_1518(dataOut[1518]),
.io_dataOut_1519(dataOut[1519]),
.io_dataOut_1520(dataOut[1520]),
.io_dataOut_1521(dataOut[1521]),
.io_dataOut_1522(dataOut[1522]),
.io_dataOut_1523(dataOut[1523]),
.io_dataOut_1524(dataOut[1524]),
.io_dataOut_1525(dataOut[1525]),
.io_dataOut_1526(dataOut[1526]),
.io_dataOut_1527(dataOut[1527]),
.io_dataOut_1528(dataOut[1528]),
.io_dataOut_1529(dataOut[1529]),
.io_dataOut_1530(dataOut[1530]),
.io_dataOut_1531(dataOut[1531]),
.io_dataOut_1532(dataOut[1532]),
.io_dataOut_1533(dataOut[1533]),
.io_dataOut_1534(dataOut[1534]),
.io_dataOut_1535(dataOut[1535]),
.io_dataOut_1536(dataOut[1536]),
.io_dataOut_1537(dataOut[1537]),
.io_dataOut_1538(dataOut[1538]),
.io_dataOut_1539(dataOut[1539]),
.io_dataOut_1540(dataOut[1540]),
.io_dataOut_1541(dataOut[1541]),
.io_dataOut_1542(dataOut[1542]),
.io_dataOut_1543(dataOut[1543]),
.io_dataOut_1544(dataOut[1544]),
.io_dataOut_1545(dataOut[1545]),
.io_dataOut_1546(dataOut[1546]),
.io_dataOut_1547(dataOut[1547]),
.io_dataOut_1548(dataOut[1548]),
.io_dataOut_1549(dataOut[1549]),
.io_dataOut_1550(dataOut[1550]),
.io_dataOut_1551(dataOut[1551]),
.io_dataOut_1552(dataOut[1552]),
.io_dataOut_1553(dataOut[1553]),
.io_dataOut_1554(dataOut[1554]),
.io_dataOut_1555(dataOut[1555]),
.io_dataOut_1556(dataOut[1556]),
.io_dataOut_1557(dataOut[1557]),
.io_dataOut_1558(dataOut[1558]),
.io_dataOut_1559(dataOut[1559]),
.io_dataOut_1560(dataOut[1560]),
.io_dataOut_1561(dataOut[1561]),
.io_dataOut_1562(dataOut[1562]),
.io_dataOut_1563(dataOut[1563]),
.io_dataOut_1564(dataOut[1564]),
.io_dataOut_1565(dataOut[1565]),
.io_dataOut_1566(dataOut[1566]),
.io_dataOut_1567(dataOut[1567]),
.io_dataOut_1568(dataOut[1568]),
.io_dataOut_1569(dataOut[1569]),
.io_dataOut_1570(dataOut[1570]),
.io_dataOut_1571(dataOut[1571]),
.io_dataOut_1572(dataOut[1572]),
.io_dataOut_1573(dataOut[1573]),
.io_dataOut_1574(dataOut[1574]),
.io_dataOut_1575(dataOut[1575]),
.io_dataOut_1576(dataOut[1576]),
.io_dataOut_1577(dataOut[1577]),
.io_dataOut_1578(dataOut[1578]),
.io_dataOut_1579(dataOut[1579]),
.io_dataOut_1580(dataOut[1580]),
.io_dataOut_1581(dataOut[1581]),
.io_dataOut_1582(dataOut[1582]),
.io_dataOut_1583(dataOut[1583]),
.io_dataOut_1584(dataOut[1584]),
.io_dataOut_1585(dataOut[1585]),
.io_dataOut_1586(dataOut[1586]),
.io_dataOut_1587(dataOut[1587]),
.io_dataOut_1588(dataOut[1588]),
.io_dataOut_1589(dataOut[1589]),
.io_dataOut_1590(dataOut[1590]),
.io_dataOut_1591(dataOut[1591]),
.io_dataOut_1592(dataOut[1592]),
.io_dataOut_1593(dataOut[1593]),
.io_dataOut_1594(dataOut[1594]),
.io_dataOut_1595(dataOut[1595]),
.io_dataOut_1596(dataOut[1596]),
.io_dataOut_1597(dataOut[1597]),
.io_dataOut_1598(dataOut[1598]),
.io_dataOut_1599(dataOut[1599]),
.io_dataOut_1600(dataOut[1600]),
.io_dataOut_1601(dataOut[1601]),
.io_dataOut_1602(dataOut[1602]),
.io_dataOut_1603(dataOut[1603]),
.io_dataOut_1604(dataOut[1604]),
.io_dataOut_1605(dataOut[1605]),
.io_dataOut_1606(dataOut[1606]),
.io_dataOut_1607(dataOut[1607]),
.io_dataOut_1608(dataOut[1608]),
.io_dataOut_1609(dataOut[1609]),
.io_dataOut_1610(dataOut[1610]),
.io_dataOut_1611(dataOut[1611]),
.io_dataOut_1612(dataOut[1612]),
.io_dataOut_1613(dataOut[1613]),
.io_dataOut_1614(dataOut[1614]),
.io_dataOut_1615(dataOut[1615]),
.io_dataOut_1616(dataOut[1616]),
.io_dataOut_1617(dataOut[1617]),
.io_dataOut_1618(dataOut[1618]),
.io_dataOut_1619(dataOut[1619]),
.io_dataOut_1620(dataOut[1620]),
.io_dataOut_1621(dataOut[1621]),
.io_dataOut_1622(dataOut[1622]),
.io_dataOut_1623(dataOut[1623]),
.io_dataOut_1624(dataOut[1624]),
.io_dataOut_1625(dataOut[1625]),
.io_dataOut_1626(dataOut[1626]),
.io_dataOut_1627(dataOut[1627]),
.io_dataOut_1628(dataOut[1628]),
.io_dataOut_1629(dataOut[1629]),
.io_dataOut_1630(dataOut[1630]),
.io_dataOut_1631(dataOut[1631]),
.io_dataOut_1632(dataOut[1632]),
.io_dataOut_1633(dataOut[1633]),
.io_dataOut_1634(dataOut[1634]),
.io_dataOut_1635(dataOut[1635]),
.io_dataOut_1636(dataOut[1636]),
.io_dataOut_1637(dataOut[1637]),
.io_dataOut_1638(dataOut[1638]),
.io_dataOut_1639(dataOut[1639]),
.io_dataOut_1640(dataOut[1640]),
.io_dataOut_1641(dataOut[1641]),
.io_dataOut_1642(dataOut[1642]),
.io_dataOut_1643(dataOut[1643]),
.io_dataOut_1644(dataOut[1644]),
.io_dataOut_1645(dataOut[1645]),
.io_dataOut_1646(dataOut[1646]),
.io_dataOut_1647(dataOut[1647]),
.io_dataOut_1648(dataOut[1648]),
.io_dataOut_1649(dataOut[1649]),
.io_dataOut_1650(dataOut[1650]),
.io_dataOut_1651(dataOut[1651]),
.io_dataOut_1652(dataOut[1652]),
.io_dataOut_1653(dataOut[1653]),
.io_dataOut_1654(dataOut[1654]),
.io_dataOut_1655(dataOut[1655]),
.io_dataOut_1656(dataOut[1656]),
.io_dataOut_1657(dataOut[1657]),
.io_dataOut_1658(dataOut[1658]),
.io_dataOut_1659(dataOut[1659]),
.io_dataOut_1660(dataOut[1660]),
.io_dataOut_1661(dataOut[1661]),
.io_dataOut_1662(dataOut[1662]),
.io_dataOut_1663(dataOut[1663]),
.io_dataOut_1664(dataOut[1664]),
.io_dataOut_1665(dataOut[1665]),
.io_dataOut_1666(dataOut[1666]),
.io_dataOut_1667(dataOut[1667]),
.io_dataOut_1668(dataOut[1668]),
.io_dataOut_1669(dataOut[1669]),
.io_dataOut_1670(dataOut[1670]),
.io_dataOut_1671(dataOut[1671]),
.io_dataOut_1672(dataOut[1672]),
.io_dataOut_1673(dataOut[1673]),
.io_dataOut_1674(dataOut[1674]),
.io_dataOut_1675(dataOut[1675]),
.io_dataOut_1676(dataOut[1676]),
.io_dataOut_1677(dataOut[1677]),
.io_dataOut_1678(dataOut[1678]),
.io_dataOut_1679(dataOut[1679]),
.io_dataOut_1680(dataOut[1680]),
.io_dataOut_1681(dataOut[1681]),
.io_dataOut_1682(dataOut[1682]),
.io_dataOut_1683(dataOut[1683]),
.io_dataOut_1684(dataOut[1684]),
.io_dataOut_1685(dataOut[1685]),
.io_dataOut_1686(dataOut[1686]),
.io_dataOut_1687(dataOut[1687]),
.io_dataOut_1688(dataOut[1688]),
.io_dataOut_1689(dataOut[1689]),
.io_dataOut_1690(dataOut[1690]),
.io_dataOut_1691(dataOut[1691]),
.io_dataOut_1692(dataOut[1692]),
.io_dataOut_1693(dataOut[1693]),
.io_dataOut_1694(dataOut[1694]),
.io_dataOut_1695(dataOut[1695]),
.io_dataOut_1696(dataOut[1696]),
.io_dataOut_1697(dataOut[1697]),
.io_dataOut_1698(dataOut[1698]),
.io_dataOut_1699(dataOut[1699]),
.io_dataOut_1700(dataOut[1700]),
.io_dataOut_1701(dataOut[1701]),
.io_dataOut_1702(dataOut[1702]),
.io_dataOut_1703(dataOut[1703]),
.io_dataOut_1704(dataOut[1704]),
.io_dataOut_1705(dataOut[1705]),
.io_dataOut_1706(dataOut[1706]),
.io_dataOut_1707(dataOut[1707]),
.io_dataOut_1708(dataOut[1708]),
.io_dataOut_1709(dataOut[1709]),
.io_dataOut_1710(dataOut[1710]),
.io_dataOut_1711(dataOut[1711]),
.io_dataOut_1712(dataOut[1712]),
.io_dataOut_1713(dataOut[1713]),
.io_dataOut_1714(dataOut[1714]),
.io_dataOut_1715(dataOut[1715]),
.io_dataOut_1716(dataOut[1716]),
.io_dataOut_1717(dataOut[1717]),
.io_dataOut_1718(dataOut[1718]),
.io_dataOut_1719(dataOut[1719]),
.io_dataOut_1720(dataOut[1720]),
.io_dataOut_1721(dataOut[1721]),
.io_dataOut_1722(dataOut[1722]),
.io_dataOut_1723(dataOut[1723]),
.io_dataOut_1724(dataOut[1724]),
.io_dataOut_1725(dataOut[1725]),
.io_dataOut_1726(dataOut[1726]),
.io_dataOut_1727(dataOut[1727]),
.io_dataOut_1728(dataOut[1728]),
.io_dataOut_1729(dataOut[1729]),
.io_dataOut_1730(dataOut[1730]),
.io_dataOut_1731(dataOut[1731]),
.io_dataOut_1732(dataOut[1732]),
.io_dataOut_1733(dataOut[1733]),
.io_dataOut_1734(dataOut[1734]),
.io_dataOut_1735(dataOut[1735]),
.io_dataOut_1736(dataOut[1736]),
.io_dataOut_1737(dataOut[1737]),
.io_dataOut_1738(dataOut[1738]),
.io_dataOut_1739(dataOut[1739]),
.io_dataOut_1740(dataOut[1740]),
.io_dataOut_1741(dataOut[1741]),
.io_dataOut_1742(dataOut[1742]),
.io_dataOut_1743(dataOut[1743]),
.io_dataOut_1744(dataOut[1744]),
.io_dataOut_1745(dataOut[1745]),
.io_dataOut_1746(dataOut[1746]),
.io_dataOut_1747(dataOut[1747]),
.io_dataOut_1748(dataOut[1748]),
.io_dataOut_1749(dataOut[1749]),
.io_dataOut_1750(dataOut[1750]),
.io_dataOut_1751(dataOut[1751]),
.io_dataOut_1752(dataOut[1752]),
.io_dataOut_1753(dataOut[1753]),
.io_dataOut_1754(dataOut[1754]),
.io_dataOut_1755(dataOut[1755]),
.io_dataOut_1756(dataOut[1756]),
.io_dataOut_1757(dataOut[1757]),
.io_dataOut_1758(dataOut[1758]),
.io_dataOut_1759(dataOut[1759]),
.io_dataOut_1760(dataOut[1760]),
.io_dataOut_1761(dataOut[1761]),
.io_dataOut_1762(dataOut[1762]),
.io_dataOut_1763(dataOut[1763]),
.io_dataOut_1764(dataOut[1764]),
.io_dataOut_1765(dataOut[1765]),
.io_dataOut_1766(dataOut[1766]),
.io_dataOut_1767(dataOut[1767]),
.io_dataOut_1768(dataOut[1768]),
.io_dataOut_1769(dataOut[1769]),
.io_dataOut_1770(dataOut[1770]),
.io_dataOut_1771(dataOut[1771]),
.io_dataOut_1772(dataOut[1772]),
.io_dataOut_1773(dataOut[1773]),
.io_dataOut_1774(dataOut[1774]),
.io_dataOut_1775(dataOut[1775]),
.io_dataOut_1776(dataOut[1776]),
.io_dataOut_1777(dataOut[1777]),
.io_dataOut_1778(dataOut[1778]),
.io_dataOut_1779(dataOut[1779]),
.io_dataOut_1780(dataOut[1780]),
.io_dataOut_1781(dataOut[1781]),
.io_dataOut_1782(dataOut[1782]),
.io_dataOut_1783(dataOut[1783]),
.io_dataOut_1784(dataOut[1784]),
.io_dataOut_1785(dataOut[1785]),
.io_dataOut_1786(dataOut[1786]),
.io_dataOut_1787(dataOut[1787]),
.io_dataOut_1788(dataOut[1788]),
.io_dataOut_1789(dataOut[1789]),
.io_dataOut_1790(dataOut[1790]),
.io_dataOut_1791(dataOut[1791]),
.io_dataOut_1792(dataOut[1792]),
.io_dataOut_1793(dataOut[1793]),
.io_dataOut_1794(dataOut[1794]),
.io_dataOut_1795(dataOut[1795]),
.io_dataOut_1796(dataOut[1796]),
.io_dataOut_1797(dataOut[1797]),
.io_dataOut_1798(dataOut[1798]),
.io_dataOut_1799(dataOut[1799]),
.io_dataOut_1800(dataOut[1800]),
.io_dataOut_1801(dataOut[1801]),
.io_dataOut_1802(dataOut[1802]),
.io_dataOut_1803(dataOut[1803]),
.io_dataOut_1804(dataOut[1804]),
.io_dataOut_1805(dataOut[1805]),
.io_dataOut_1806(dataOut[1806]),
.io_dataOut_1807(dataOut[1807]),
.io_dataOut_1808(dataOut[1808]),
.io_dataOut_1809(dataOut[1809]),
.io_dataOut_1810(dataOut[1810]),
.io_dataOut_1811(dataOut[1811]),
.io_dataOut_1812(dataOut[1812]),
.io_dataOut_1813(dataOut[1813]),
.io_dataOut_1814(dataOut[1814]),
.io_dataOut_1815(dataOut[1815]),
.io_dataOut_1816(dataOut[1816]),
.io_dataOut_1817(dataOut[1817]),
.io_dataOut_1818(dataOut[1818]),
.io_dataOut_1819(dataOut[1819]),
.io_dataOut_1820(dataOut[1820]),
.io_dataOut_1821(dataOut[1821]),
.io_dataOut_1822(dataOut[1822]),
.io_dataOut_1823(dataOut[1823]),
.io_dataOut_1824(dataOut[1824]),
.io_dataOut_1825(dataOut[1825]),
.io_dataOut_1826(dataOut[1826]),
.io_dataOut_1827(dataOut[1827]),
.io_dataOut_1828(dataOut[1828]),
.io_dataOut_1829(dataOut[1829]),
.io_dataOut_1830(dataOut[1830]),
.io_dataOut_1831(dataOut[1831]),
.io_dataOut_1832(dataOut[1832]),
.io_dataOut_1833(dataOut[1833]),
.io_dataOut_1834(dataOut[1834]),
.io_dataOut_1835(dataOut[1835]),
.io_dataOut_1836(dataOut[1836]),
.io_dataOut_1837(dataOut[1837]),
.io_dataOut_1838(dataOut[1838]),
.io_dataOut_1839(dataOut[1839]),
.io_dataOut_1840(dataOut[1840]),
.io_dataOut_1841(dataOut[1841]),
.io_dataOut_1842(dataOut[1842]),
.io_dataOut_1843(dataOut[1843]),
.io_dataOut_1844(dataOut[1844]),
.io_dataOut_1845(dataOut[1845]),
.io_dataOut_1846(dataOut[1846]),
.io_dataOut_1847(dataOut[1847]),
.io_dataOut_1848(dataOut[1848]),
.io_dataOut_1849(dataOut[1849]),
.io_dataOut_1850(dataOut[1850]),
.io_dataOut_1851(dataOut[1851]),
.io_dataOut_1852(dataOut[1852]),
.io_dataOut_1853(dataOut[1853]),
.io_dataOut_1854(dataOut[1854]),
.io_dataOut_1855(dataOut[1855]),
.io_dataOut_1856(dataOut[1856]),
.io_dataOut_1857(dataOut[1857]),
.io_dataOut_1858(dataOut[1858]),
.io_dataOut_1859(dataOut[1859]),
.io_dataOut_1860(dataOut[1860]),
.io_dataOut_1861(dataOut[1861]),
.io_dataOut_1862(dataOut[1862]),
.io_dataOut_1863(dataOut[1863]),
.io_dataOut_1864(dataOut[1864]),
.io_dataOut_1865(dataOut[1865]),
.io_dataOut_1866(dataOut[1866]),
.io_dataOut_1867(dataOut[1867]),
.io_dataOut_1868(dataOut[1868]),
.io_dataOut_1869(dataOut[1869]),
.io_dataOut_1870(dataOut[1870]),
.io_dataOut_1871(dataOut[1871]),
.io_dataOut_1872(dataOut[1872]),
.io_dataOut_1873(dataOut[1873]),
.io_dataOut_1874(dataOut[1874]),
.io_dataOut_1875(dataOut[1875]),
.io_dataOut_1876(dataOut[1876]),
.io_dataOut_1877(dataOut[1877]),
.io_dataOut_1878(dataOut[1878]),
.io_dataOut_1879(dataOut[1879]),
.io_dataOut_1880(dataOut[1880]),
.io_dataOut_1881(dataOut[1881]),
.io_dataOut_1882(dataOut[1882]),
.io_dataOut_1883(dataOut[1883]),
.io_dataOut_1884(dataOut[1884]),
.io_dataOut_1885(dataOut[1885]),
.io_dataOut_1886(dataOut[1886]),
.io_dataOut_1887(dataOut[1887]),
.io_dataOut_1888(dataOut[1888]),
.io_dataOut_1889(dataOut[1889]),
.io_dataOut_1890(dataOut[1890]),
.io_dataOut_1891(dataOut[1891]),
.io_dataOut_1892(dataOut[1892]),
.io_dataOut_1893(dataOut[1893]),
.io_dataOut_1894(dataOut[1894]),
.io_dataOut_1895(dataOut[1895]),
.io_dataOut_1896(dataOut[1896]),
.io_dataOut_1897(dataOut[1897]),
.io_dataOut_1898(dataOut[1898]),
.io_dataOut_1899(dataOut[1899]),
.io_dataOut_1900(dataOut[1900]),
.io_dataOut_1901(dataOut[1901]),
.io_dataOut_1902(dataOut[1902]),
.io_dataOut_1903(dataOut[1903]),
.io_dataOut_1904(dataOut[1904]),
.io_dataOut_1905(dataOut[1905]),
.io_dataOut_1906(dataOut[1906]),
.io_dataOut_1907(dataOut[1907]),
.io_dataOut_1908(dataOut[1908]),
.io_dataOut_1909(dataOut[1909]),
.io_dataOut_1910(dataOut[1910]),
.io_dataOut_1911(dataOut[1911]),
.io_dataOut_1912(dataOut[1912]),
.io_dataOut_1913(dataOut[1913]),
.io_dataOut_1914(dataOut[1914]),
.io_dataOut_1915(dataOut[1915]),
.io_dataOut_1916(dataOut[1916]),
.io_dataOut_1917(dataOut[1917]),
.io_dataOut_1918(dataOut[1918]),
.io_dataOut_1919(dataOut[1919]),
.io_dataOut_1920(dataOut[1920]),
.io_dataOut_1921(dataOut[1921]),
.io_dataOut_1922(dataOut[1922]),
.io_dataOut_1923(dataOut[1923]),
.io_dataOut_1924(dataOut[1924]),
.io_dataOut_1925(dataOut[1925]),
.io_dataOut_1926(dataOut[1926]),
.io_dataOut_1927(dataOut[1927]),
.io_dataOut_1928(dataOut[1928]),
.io_dataOut_1929(dataOut[1929]),
.io_dataOut_1930(dataOut[1930]),
.io_dataOut_1931(dataOut[1931]),
.io_dataOut_1932(dataOut[1932]),
.io_dataOut_1933(dataOut[1933]),
.io_dataOut_1934(dataOut[1934]),
.io_dataOut_1935(dataOut[1935]),
.io_dataOut_1936(dataOut[1936]),
.io_dataOut_1937(dataOut[1937]),
.io_dataOut_1938(dataOut[1938]),
.io_dataOut_1939(dataOut[1939]),
.io_dataOut_1940(dataOut[1940]),
.io_dataOut_1941(dataOut[1941]),
.io_dataOut_1942(dataOut[1942]),
.io_dataOut_1943(dataOut[1943]),
.io_dataOut_1944(dataOut[1944]),
.io_dataOut_1945(dataOut[1945]),
.io_dataOut_1946(dataOut[1946]),
.io_dataOut_1947(dataOut[1947]),
.io_dataOut_1948(dataOut[1948]),
.io_dataOut_1949(dataOut[1949]),
.io_dataOut_1950(dataOut[1950]),
.io_dataOut_1951(dataOut[1951]),
.io_dataOut_1952(dataOut[1952]),
.io_dataOut_1953(dataOut[1953]),
.io_dataOut_1954(dataOut[1954]),
.io_dataOut_1955(dataOut[1955]),
.io_dataOut_1956(dataOut[1956]),
.io_dataOut_1957(dataOut[1957]),
.io_dataOut_1958(dataOut[1958]),
.io_dataOut_1959(dataOut[1959]),
.io_dataOut_1960(dataOut[1960]),
.io_dataOut_1961(dataOut[1961]),
.io_dataOut_1962(dataOut[1962]),
.io_dataOut_1963(dataOut[1963]),
.io_dataOut_1964(dataOut[1964]),
.io_dataOut_1965(dataOut[1965]),
.io_dataOut_1966(dataOut[1966]),
.io_dataOut_1967(dataOut[1967]),
.io_dataOut_1968(dataOut[1968]),
.io_dataOut_1969(dataOut[1969]),
.io_dataOut_1970(dataOut[1970]),
.io_dataOut_1971(dataOut[1971]),
.io_dataOut_1972(dataOut[1972]),
.io_dataOut_1973(dataOut[1973]),
.io_dataOut_1974(dataOut[1974]),
.io_dataOut_1975(dataOut[1975]),
.io_dataOut_1976(dataOut[1976]),
.io_dataOut_1977(dataOut[1977]),
.io_dataOut_1978(dataOut[1978]),
.io_dataOut_1979(dataOut[1979]),
.io_dataOut_1980(dataOut[1980]),
.io_dataOut_1981(dataOut[1981]),
.io_dataOut_1982(dataOut[1982]),
.io_dataOut_1983(dataOut[1983]),
.io_dataOut_1984(dataOut[1984]),
.io_dataOut_1985(dataOut[1985]),
.io_dataOut_1986(dataOut[1986]),
.io_dataOut_1987(dataOut[1987]),
.io_dataOut_1988(dataOut[1988]),
.io_dataOut_1989(dataOut[1989]),
.io_dataOut_1990(dataOut[1990]),
.io_dataOut_1991(dataOut[1991]),
.io_dataOut_1992(dataOut[1992]),
.io_dataOut_1993(dataOut[1993]),
.io_dataOut_1994(dataOut[1994]),
.io_dataOut_1995(dataOut[1995]),
.io_dataOut_1996(dataOut[1996]),
.io_dataOut_1997(dataOut[1997]),
.io_dataOut_1998(dataOut[1998]),
.io_dataOut_1999(dataOut[1999]),
.io_dataOut_2000(dataOut[2000]),
.io_dataOut_2001(dataOut[2001]),
.io_dataOut_2002(dataOut[2002]),
.io_dataOut_2003(dataOut[2003]),
.io_dataOut_2004(dataOut[2004]),
.io_dataOut_2005(dataOut[2005]),
.io_dataOut_2006(dataOut[2006]),
.io_dataOut_2007(dataOut[2007]),
.io_dataOut_2008(dataOut[2008]),
.io_dataOut_2009(dataOut[2009]),
.io_dataOut_2010(dataOut[2010]),
.io_dataOut_2011(dataOut[2011]),
.io_dataOut_2012(dataOut[2012]),
.io_dataOut_2013(dataOut[2013]),
.io_dataOut_2014(dataOut[2014]),
.io_dataOut_2015(dataOut[2015]),
.io_dataOut_2016(dataOut[2016]),
.io_dataOut_2017(dataOut[2017]),
.io_dataOut_2018(dataOut[2018]),
.io_dataOut_2019(dataOut[2019]),
.io_dataOut_2020(dataOut[2020]),
.io_dataOut_2021(dataOut[2021]),
.io_dataOut_2022(dataOut[2022]),
.io_dataOut_2023(dataOut[2023]),
.io_dataOut_2024(dataOut[2024]),
.io_dataOut_2025(dataOut[2025]),
.io_dataOut_2026(dataOut[2026]),
.io_dataOut_2027(dataOut[2027]),
.io_dataOut_2028(dataOut[2028]),
.io_dataOut_2029(dataOut[2029]),
.io_dataOut_2030(dataOut[2030]),
.io_dataOut_2031(dataOut[2031]),
.io_dataOut_2032(dataOut[2032]),
.io_dataOut_2033(dataOut[2033]),
.io_dataOut_2034(dataOut[2034]),
.io_dataOut_2035(dataOut[2035]),
.io_dataOut_2036(dataOut[2036]),
.io_dataOut_2037(dataOut[2037]),
.io_dataOut_2038(dataOut[2038]),
.io_dataOut_2039(dataOut[2039]),
.io_dataOut_2040(dataOut[2040]),
.io_dataOut_2041(dataOut[2041]),
.io_dataOut_2042(dataOut[2042]),
.io_dataOut_2043(dataOut[2043]),
.io_dataOut_2044(dataOut[2044]),
.io_dataOut_2045(dataOut[2045]),
.io_dataOut_2046(dataOut[2046]),
.io_dataOut_2047(dataOut[2047]),
.io_dataOut_2048(dataOut[2048]),
.io_dataOut_2049(dataOut[2049]),
.io_dataOut_2050(dataOut[2050]),
.io_dataOut_2051(dataOut[2051]),
.io_dataOut_2052(dataOut[2052]),
.io_dataOut_2053(dataOut[2053]),
.io_dataOut_2054(dataOut[2054]),
.io_dataOut_2055(dataOut[2055]),
.io_dataOut_2056(dataOut[2056]),
.io_dataOut_2057(dataOut[2057]),
.io_dataOut_2058(dataOut[2058]),
.io_dataOut_2059(dataOut[2059]),
.io_dataOut_2060(dataOut[2060]),
.io_dataOut_2061(dataOut[2061]),
.io_dataOut_2062(dataOut[2062]),
.io_dataOut_2063(dataOut[2063]),
.io_dataOut_2064(dataOut[2064]),
.io_dataOut_2065(dataOut[2065]),
.io_dataOut_2066(dataOut[2066]),
.io_dataOut_2067(dataOut[2067]),
.io_dataOut_2068(dataOut[2068]),
.io_dataOut_2069(dataOut[2069]),
.io_dataOut_2070(dataOut[2070]),
.io_dataOut_2071(dataOut[2071]),
.io_dataOut_2072(dataOut[2072]),
.io_dataOut_2073(dataOut[2073]),
.io_dataOut_2074(dataOut[2074]),
.io_dataOut_2075(dataOut[2075]),
.io_dataOut_2076(dataOut[2076]),
.io_dataOut_2077(dataOut[2077]),
.io_dataOut_2078(dataOut[2078]),
.io_dataOut_2079(dataOut[2079]),
.io_dataOut_2080(dataOut[2080]),
.io_dataOut_2081(dataOut[2081]),
.io_dataOut_2082(dataOut[2082]),
.io_dataOut_2083(dataOut[2083]),
.io_dataOut_2084(dataOut[2084]),
.io_dataOut_2085(dataOut[2085]),
.io_dataOut_2086(dataOut[2086]),
.io_dataOut_2087(dataOut[2087]),
.io_dataOut_2088(dataOut[2088]),
.io_dataOut_2089(dataOut[2089]),
.io_dataOut_2090(dataOut[2090]),
.io_dataOut_2091(dataOut[2091]),
.io_dataOut_2092(dataOut[2092]),
.io_dataOut_2093(dataOut[2093]),
.io_dataOut_2094(dataOut[2094]),
.io_dataOut_2095(dataOut[2095]),
.io_dataOut_2096(dataOut[2096]),
.io_dataOut_2097(dataOut[2097]),
.io_dataOut_2098(dataOut[2098]),
.io_dataOut_2099(dataOut[2099]),
.io_dataOut_2100(dataOut[2100]),
.io_dataOut_2101(dataOut[2101]),
.io_dataOut_2102(dataOut[2102]),
.io_dataOut_2103(dataOut[2103]),
.io_dataOut_2104(dataOut[2104]),
.io_dataOut_2105(dataOut[2105]),
.io_dataOut_2106(dataOut[2106]),
.io_dataOut_2107(dataOut[2107]),
.io_dataOut_2108(dataOut[2108]),
.io_dataOut_2109(dataOut[2109]),
.io_dataOut_2110(dataOut[2110]),
.io_dataOut_2111(dataOut[2111]),
.io_dataOut_2112(dataOut[2112]),
.io_dataOut_2113(dataOut[2113]),
.io_dataOut_2114(dataOut[2114]),
.io_dataOut_2115(dataOut[2115]),
.io_dataOut_2116(dataOut[2116]),
.io_dataOut_2117(dataOut[2117]),
.io_dataOut_2118(dataOut[2118]),
.io_dataOut_2119(dataOut[2119]),
.io_dataOut_2120(dataOut[2120]),
.io_dataOut_2121(dataOut[2121]),
.io_dataOut_2122(dataOut[2122]),
.io_dataOut_2123(dataOut[2123]),
.io_dataOut_2124(dataOut[2124]),
.io_dataOut_2125(dataOut[2125]),
.io_dataOut_2126(dataOut[2126]),
.io_dataOut_2127(dataOut[2127]),
.io_dataOut_2128(dataOut[2128]),
.io_dataOut_2129(dataOut[2129]),
.io_dataOut_2130(dataOut[2130]),
.io_dataOut_2131(dataOut[2131]),
.io_dataOut_2132(dataOut[2132]),
.io_dataOut_2133(dataOut[2133]),
.io_dataOut_2134(dataOut[2134]),
.io_dataOut_2135(dataOut[2135]),
.io_dataOut_2136(dataOut[2136]),
.io_dataOut_2137(dataOut[2137]),
.io_dataOut_2138(dataOut[2138]),
.io_dataOut_2139(dataOut[2139]),
.io_dataOut_2140(dataOut[2140]),
.io_dataOut_2141(dataOut[2141]),
.io_dataOut_2142(dataOut[2142]),
.io_dataOut_2143(dataOut[2143]),
.io_dataOut_2144(dataOut[2144]),
.io_dataOut_2145(dataOut[2145]),
.io_dataOut_2146(dataOut[2146]),
.io_dataOut_2147(dataOut[2147]),
.io_dataOut_2148(dataOut[2148]),
.io_dataOut_2149(dataOut[2149]),
.io_dataOut_2150(dataOut[2150]),
.io_dataOut_2151(dataOut[2151]),
.io_dataOut_2152(dataOut[2152]),
.io_dataOut_2153(dataOut[2153]),
.io_dataOut_2154(dataOut[2154]),
.io_dataOut_2155(dataOut[2155]),
.io_dataOut_2156(dataOut[2156]),
.io_dataOut_2157(dataOut[2157]),
.io_dataOut_2158(dataOut[2158]),
.io_dataOut_2159(dataOut[2159]),
.io_dataOut_2160(dataOut[2160]),
.io_dataOut_2161(dataOut[2161]),
.io_dataOut_2162(dataOut[2162]),
.io_dataOut_2163(dataOut[2163]),
.io_dataOut_2164(dataOut[2164]),
.io_dataOut_2165(dataOut[2165]),
.io_dataOut_2166(dataOut[2166]),
.io_dataOut_2167(dataOut[2167]),
.io_dataOut_2168(dataOut[2168]),
.io_dataOut_2169(dataOut[2169]),
.io_dataOut_2170(dataOut[2170]),
.io_dataOut_2171(dataOut[2171]),
.io_dataOut_2172(dataOut[2172]),
.io_dataOut_2173(dataOut[2173]),
.io_dataOut_2174(dataOut[2174]),
.io_dataOut_2175(dataOut[2175]),
.io_dataOut_2176(dataOut[2176]),
.io_dataOut_2177(dataOut[2177]),
.io_dataOut_2178(dataOut[2178]),
.io_dataOut_2179(dataOut[2179]),
.io_dataOut_2180(dataOut[2180]),
.io_dataOut_2181(dataOut[2181]),
.io_dataOut_2182(dataOut[2182]),
.io_dataOut_2183(dataOut[2183]),
.io_dataOut_2184(dataOut[2184]),
.io_dataOut_2185(dataOut[2185]),
.io_dataOut_2186(dataOut[2186]),
.io_dataOut_2187(dataOut[2187]),
.io_dataOut_2188(dataOut[2188]),
.io_dataOut_2189(dataOut[2189]),
.io_dataOut_2190(dataOut[2190]),
.io_dataOut_2191(dataOut[2191]),
.io_dataOut_2192(dataOut[2192]),
.io_dataOut_2193(dataOut[2193]),
.io_dataOut_2194(dataOut[2194]),
.io_dataOut_2195(dataOut[2195]),
.io_dataOut_2196(dataOut[2196]),
.io_dataOut_2197(dataOut[2197]),
.io_dataOut_2198(dataOut[2198]),
.io_dataOut_2199(dataOut[2199]),
.io_dataOut_2200(dataOut[2200]),
.io_dataOut_2201(dataOut[2201]),
.io_dataOut_2202(dataOut[2202]),
.io_dataOut_2203(dataOut[2203]),
.io_dataOut_2204(dataOut[2204]),
.io_dataOut_2205(dataOut[2205]),
.io_dataOut_2206(dataOut[2206]),
.io_dataOut_2207(dataOut[2207]),
.io_dataOut_2208(dataOut[2208]),
.io_dataOut_2209(dataOut[2209]),
.io_dataOut_2210(dataOut[2210]),
.io_dataOut_2211(dataOut[2211]),
.io_dataOut_2212(dataOut[2212]),
.io_dataOut_2213(dataOut[2213]),
.io_dataOut_2214(dataOut[2214]),
.io_dataOut_2215(dataOut[2215]),
.io_dataOut_2216(dataOut[2216]),
.io_dataOut_2217(dataOut[2217]),
.io_dataOut_2218(dataOut[2218]),
.io_dataOut_2219(dataOut[2219]),
.io_dataOut_2220(dataOut[2220]),
.io_dataOut_2221(dataOut[2221]),
.io_dataOut_2222(dataOut[2222]),
.io_dataOut_2223(dataOut[2223]),
.io_dataOut_2224(dataOut[2224]),
.io_dataOut_2225(dataOut[2225]),
.io_dataOut_2226(dataOut[2226]),
.io_dataOut_2227(dataOut[2227]),
.io_dataOut_2228(dataOut[2228]),
.io_dataOut_2229(dataOut[2229]),
.io_dataOut_2230(dataOut[2230]),
.io_dataOut_2231(dataOut[2231]),
.io_dataOut_2232(dataOut[2232]),
.io_dataOut_2233(dataOut[2233]),
.io_dataOut_2234(dataOut[2234]),
.io_dataOut_2235(dataOut[2235]),
.io_dataOut_2236(dataOut[2236]),
.io_dataOut_2237(dataOut[2237]),
.io_dataOut_2238(dataOut[2238]),
.io_dataOut_2239(dataOut[2239]),
.io_dataOut_2240(dataOut[2240]),
.io_dataOut_2241(dataOut[2241]),
.io_dataOut_2242(dataOut[2242]),
.io_dataOut_2243(dataOut[2243]),
.io_dataOut_2244(dataOut[2244]),
.io_dataOut_2245(dataOut[2245]),
.io_dataOut_2246(dataOut[2246]),
.io_dataOut_2247(dataOut[2247]),
.io_dataOut_2248(dataOut[2248]),
.io_dataOut_2249(dataOut[2249]),
.io_dataOut_2250(dataOut[2250]),
.io_dataOut_2251(dataOut[2251]),
.io_dataOut_2252(dataOut[2252]),
.io_dataOut_2253(dataOut[2253]),
.io_dataOut_2254(dataOut[2254]),
.io_dataOut_2255(dataOut[2255]),
.io_dataOut_2256(dataOut[2256]),
.io_dataOut_2257(dataOut[2257]),
.io_dataOut_2258(dataOut[2258]),
.io_dataOut_2259(dataOut[2259]),
.io_dataOut_2260(dataOut[2260]),
.io_dataOut_2261(dataOut[2261]),
.io_dataOut_2262(dataOut[2262]),
.io_dataOut_2263(dataOut[2263]),
.io_dataOut_2264(dataOut[2264]),
.io_dataOut_2265(dataOut[2265]),
.io_dataOut_2266(dataOut[2266]),
.io_dataOut_2267(dataOut[2267]),
.io_dataOut_2268(dataOut[2268]),
.io_dataOut_2269(dataOut[2269]),
.io_dataOut_2270(dataOut[2270]),
.io_dataOut_2271(dataOut[2271]),
.io_dataOut_2272(dataOut[2272]),
.io_dataOut_2273(dataOut[2273]),
.io_dataOut_2274(dataOut[2274]),
.io_dataOut_2275(dataOut[2275]),
.io_dataOut_2276(dataOut[2276]),
.io_dataOut_2277(dataOut[2277]),
.io_dataOut_2278(dataOut[2278]),
.io_dataOut_2279(dataOut[2279]),
.io_dataOut_2280(dataOut[2280]),
.io_dataOut_2281(dataOut[2281]),
.io_dataOut_2282(dataOut[2282]),
.io_dataOut_2283(dataOut[2283]),
.io_dataOut_2284(dataOut[2284]),
.io_dataOut_2285(dataOut[2285]),
.io_dataOut_2286(dataOut[2286]),
.io_dataOut_2287(dataOut[2287]),
.io_dataOut_2288(dataOut[2288]),
.io_dataOut_2289(dataOut[2289]),
.io_dataOut_2290(dataOut[2290]),
.io_dataOut_2291(dataOut[2291]),
.io_dataOut_2292(dataOut[2292]),
.io_dataOut_2293(dataOut[2293]),
.io_dataOut_2294(dataOut[2294]),
.io_dataOut_2295(dataOut[2295]),
.io_dataOut_2296(dataOut[2296]),
.io_dataOut_2297(dataOut[2297]),
.io_dataOut_2298(dataOut[2298]),
.io_dataOut_2299(dataOut[2299]),
.io_dataOut_2300(dataOut[2300]),
.io_dataOut_2301(dataOut[2301]),
.io_dataOut_2302(dataOut[2302]),
.io_dataOut_2303(dataOut[2303]),
.io_dataOut_2304(dataOut[2304]),
.io_dataOut_2305(dataOut[2305]),
.io_dataOut_2306(dataOut[2306]),
.io_dataOut_2307(dataOut[2307]),
.io_dataOut_2308(dataOut[2308]),
.io_dataOut_2309(dataOut[2309]),
.io_dataOut_2310(dataOut[2310]),
.io_dataOut_2311(dataOut[2311]),
.io_dataOut_2312(dataOut[2312]),
.io_dataOut_2313(dataOut[2313]),
.io_dataOut_2314(dataOut[2314]),
.io_dataOut_2315(dataOut[2315]),
.io_dataOut_2316(dataOut[2316]),
.io_dataOut_2317(dataOut[2317]),
.io_dataOut_2318(dataOut[2318]),
.io_dataOut_2319(dataOut[2319]),
.io_dataOut_2320(dataOut[2320]),
.io_dataOut_2321(dataOut[2321]),
.io_dataOut_2322(dataOut[2322]),
.io_dataOut_2323(dataOut[2323]),
.io_dataOut_2324(dataOut[2324]),
.io_dataOut_2325(dataOut[2325]),
.io_dataOut_2326(dataOut[2326]),
.io_dataOut_2327(dataOut[2327]),
.io_dataOut_2328(dataOut[2328]),
.io_dataOut_2329(dataOut[2329]),
.io_dataOut_2330(dataOut[2330]),
.io_dataOut_2331(dataOut[2331]),
.io_dataOut_2332(dataOut[2332]),
.io_dataOut_2333(dataOut[2333]),
.io_dataOut_2334(dataOut[2334]),
.io_dataOut_2335(dataOut[2335]),
.io_dataOut_2336(dataOut[2336]),
.io_dataOut_2337(dataOut[2337]),
.io_dataOut_2338(dataOut[2338]),
.io_dataOut_2339(dataOut[2339]),
.io_dataOut_2340(dataOut[2340]),
.io_dataOut_2341(dataOut[2341]),
.io_dataOut_2342(dataOut[2342]),
.io_dataOut_2343(dataOut[2343]),
.io_dataOut_2344(dataOut[2344]),
.io_dataOut_2345(dataOut[2345]),
.io_dataOut_2346(dataOut[2346]),
.io_dataOut_2347(dataOut[2347]),
.io_dataOut_2348(dataOut[2348]),
.io_dataOut_2349(dataOut[2349]),
.io_dataOut_2350(dataOut[2350]),
.io_dataOut_2351(dataOut[2351]),
.io_dataOut_2352(dataOut[2352]),
.io_dataOut_2353(dataOut[2353]),
.io_dataOut_2354(dataOut[2354]),
.io_dataOut_2355(dataOut[2355]),
.io_dataOut_2356(dataOut[2356]),
.io_dataOut_2357(dataOut[2357]),
.io_dataOut_2358(dataOut[2358]),
.io_dataOut_2359(dataOut[2359]),
.io_dataOut_2360(dataOut[2360]),
.io_dataOut_2361(dataOut[2361]),
.io_dataOut_2362(dataOut[2362]),
.io_dataOut_2363(dataOut[2363]),
.io_dataOut_2364(dataOut[2364]),
.io_dataOut_2365(dataOut[2365]),
.io_dataOut_2366(dataOut[2366]),
.io_dataOut_2367(dataOut[2367]),
.io_dataOut_2368(dataOut[2368]),
.io_dataOut_2369(dataOut[2369]),
.io_dataOut_2370(dataOut[2370]),
.io_dataOut_2371(dataOut[2371]),
.io_dataOut_2372(dataOut[2372]),
.io_dataOut_2373(dataOut[2373]),
.io_dataOut_2374(dataOut[2374]),
.io_dataOut_2375(dataOut[2375]),
.io_dataOut_2376(dataOut[2376]),
.io_dataOut_2377(dataOut[2377]),
.io_dataOut_2378(dataOut[2378]),
.io_dataOut_2379(dataOut[2379]),
.io_dataOut_2380(dataOut[2380]),
.io_dataOut_2381(dataOut[2381]),
.io_dataOut_2382(dataOut[2382]),
.io_dataOut_2383(dataOut[2383]),
.io_dataOut_2384(dataOut[2384]),
.io_dataOut_2385(dataOut[2385]),
.io_dataOut_2386(dataOut[2386]),
.io_dataOut_2387(dataOut[2387]),
.io_dataOut_2388(dataOut[2388]),
.io_dataOut_2389(dataOut[2389]),
.io_dataOut_2390(dataOut[2390]),
.io_dataOut_2391(dataOut[2391]),
.io_dataOut_2392(dataOut[2392]),
.io_dataOut_2393(dataOut[2393]),
.io_dataOut_2394(dataOut[2394]),
.io_dataOut_2395(dataOut[2395]),
.io_dataOut_2396(dataOut[2396]),
.io_dataOut_2397(dataOut[2397]),
.io_dataOut_2398(dataOut[2398]),
.io_dataOut_2399(dataOut[2399]),
.io_dataOut_2400(dataOut[2400]),
.io_dataOut_2401(dataOut[2401]),
.io_dataOut_2402(dataOut[2402]),
.io_dataOut_2403(dataOut[2403]),
.io_dataOut_2404(dataOut[2404]),
.io_dataOut_2405(dataOut[2405]),
.io_dataOut_2406(dataOut[2406]),
.io_dataOut_2407(dataOut[2407]),
.io_dataOut_2408(dataOut[2408]),
.io_dataOut_2409(dataOut[2409]),
.io_dataOut_2410(dataOut[2410]),
.io_dataOut_2411(dataOut[2411]),
.io_dataOut_2412(dataOut[2412]),
.io_dataOut_2413(dataOut[2413]),
.io_dataOut_2414(dataOut[2414]),
.io_dataOut_2415(dataOut[2415]),
.io_dataOut_2416(dataOut[2416]),
.io_dataOut_2417(dataOut[2417]),
.io_dataOut_2418(dataOut[2418]),
.io_dataOut_2419(dataOut[2419]),
.io_dataOut_2420(dataOut[2420]),
.io_dataOut_2421(dataOut[2421]),
.io_dataOut_2422(dataOut[2422]),
.io_dataOut_2423(dataOut[2423]),
.io_dataOut_2424(dataOut[2424]),
.io_dataOut_2425(dataOut[2425]),
.io_dataOut_2426(dataOut[2426]),
.io_dataOut_2427(dataOut[2427]),
.io_dataOut_2428(dataOut[2428]),
.io_dataOut_2429(dataOut[2429]),
.io_dataOut_2430(dataOut[2430]),
.io_dataOut_2431(dataOut[2431]),
.io_dataOut_2432(dataOut[2432]),
.io_dataOut_2433(dataOut[2433]),
.io_dataOut_2434(dataOut[2434]),
.io_dataOut_2435(dataOut[2435]),
.io_dataOut_2436(dataOut[2436]),
.io_dataOut_2437(dataOut[2437]),
.io_dataOut_2438(dataOut[2438]),
.io_dataOut_2439(dataOut[2439]),
.io_dataOut_2440(dataOut[2440]),
.io_dataOut_2441(dataOut[2441]),
.io_dataOut_2442(dataOut[2442]),
.io_dataOut_2443(dataOut[2443]),
.io_dataOut_2444(dataOut[2444]),
.io_dataOut_2445(dataOut[2445]),
.io_dataOut_2446(dataOut[2446]),
.io_dataOut_2447(dataOut[2447]),
.io_dataOut_2448(dataOut[2448]),
.io_dataOut_2449(dataOut[2449]),
.io_dataOut_2450(dataOut[2450]),
.io_dataOut_2451(dataOut[2451]),
.io_dataOut_2452(dataOut[2452]),
.io_dataOut_2453(dataOut[2453]),
.io_dataOut_2454(dataOut[2454]),
.io_dataOut_2455(dataOut[2455]),
.io_dataOut_2456(dataOut[2456]),
.io_dataOut_2457(dataOut[2457]),
.io_dataOut_2458(dataOut[2458]),
.io_dataOut_2459(dataOut[2459]),
.io_dataOut_2460(dataOut[2460]),
.io_dataOut_2461(dataOut[2461]),
.io_dataOut_2462(dataOut[2462]),
.io_dataOut_2463(dataOut[2463]),
.io_dataOut_2464(dataOut[2464]),
.io_dataOut_2465(dataOut[2465]),
.io_dataOut_2466(dataOut[2466]),
.io_dataOut_2467(dataOut[2467]),
.io_dataOut_2468(dataOut[2468]),
.io_dataOut_2469(dataOut[2469]),
.io_dataOut_2470(dataOut[2470]),
.io_dataOut_2471(dataOut[2471]),
.io_dataOut_2472(dataOut[2472]),
.io_dataOut_2473(dataOut[2473]),
.io_dataOut_2474(dataOut[2474]),
.io_dataOut_2475(dataOut[2475]),
.io_dataOut_2476(dataOut[2476]),
.io_dataOut_2477(dataOut[2477]),
.io_dataOut_2478(dataOut[2478]),
.io_dataOut_2479(dataOut[2479]),
.io_dataOut_2480(dataOut[2480]),
.io_dataOut_2481(dataOut[2481]),
.io_dataOut_2482(dataOut[2482]),
.io_dataOut_2483(dataOut[2483]),
.io_dataOut_2484(dataOut[2484]),
.io_dataOut_2485(dataOut[2485]),
.io_dataOut_2486(dataOut[2486]),
.io_dataOut_2487(dataOut[2487]),
.io_dataOut_2488(dataOut[2488]),
.io_dataOut_2489(dataOut[2489]),
.io_dataOut_2490(dataOut[2490]),
.io_dataOut_2491(dataOut[2491]),
.io_dataOut_2492(dataOut[2492]),
.io_dataOut_2493(dataOut[2493]),
.io_dataOut_2494(dataOut[2494]),
.io_dataOut_2495(dataOut[2495]),
.io_dataOut_2496(dataOut[2496]),
.io_dataOut_2497(dataOut[2497]),
.io_dataOut_2498(dataOut[2498]),
.io_dataOut_2499(dataOut[2499]),
.io_dataOut_2500(dataOut[2500]),
.io_dataOut_2501(dataOut[2501]),
.io_dataOut_2502(dataOut[2502]),
.io_dataOut_2503(dataOut[2503]),
.io_dataOut_2504(dataOut[2504]),
.io_dataOut_2505(dataOut[2505]),
.io_dataOut_2506(dataOut[2506]),
.io_dataOut_2507(dataOut[2507]),
.io_dataOut_2508(dataOut[2508]),
.io_dataOut_2509(dataOut[2509]),
.io_dataOut_2510(dataOut[2510]),
.io_dataOut_2511(dataOut[2511]),
.io_dataOut_2512(dataOut[2512]),
.io_dataOut_2513(dataOut[2513]),
.io_dataOut_2514(dataOut[2514]),
.io_dataOut_2515(dataOut[2515]),
.io_dataOut_2516(dataOut[2516]),
.io_dataOut_2517(dataOut[2517]),
.io_dataOut_2518(dataOut[2518]),
.io_dataOut_2519(dataOut[2519]),
.io_dataOut_2520(dataOut[2520]),
.io_dataOut_2521(dataOut[2521]),
.io_dataOut_2522(dataOut[2522]),
.io_dataOut_2523(dataOut[2523]),
.io_dataOut_2524(dataOut[2524]),
.io_dataOut_2525(dataOut[2525]),
.io_dataOut_2526(dataOut[2526]),
.io_dataOut_2527(dataOut[2527]),
.io_dataOut_2528(dataOut[2528]),
.io_dataOut_2529(dataOut[2529]),
.io_dataOut_2530(dataOut[2530]),
.io_dataOut_2531(dataOut[2531]),
.io_dataOut_2532(dataOut[2532]),
.io_dataOut_2533(dataOut[2533]),
.io_dataOut_2534(dataOut[2534]),
.io_dataOut_2535(dataOut[2535]),
.io_dataOut_2536(dataOut[2536]),
.io_dataOut_2537(dataOut[2537]),
.io_dataOut_2538(dataOut[2538]),
.io_dataOut_2539(dataOut[2539]),
.io_dataOut_2540(dataOut[2540]),
.io_dataOut_2541(dataOut[2541]),
.io_dataOut_2542(dataOut[2542]),
.io_dataOut_2543(dataOut[2543]),
.io_dataOut_2544(dataOut[2544]),
.io_dataOut_2545(dataOut[2545]),
.io_dataOut_2546(dataOut[2546]),
.io_dataOut_2547(dataOut[2547]),
.io_dataOut_2548(dataOut[2548]),
.io_dataOut_2549(dataOut[2549]),
.io_dataOut_2550(dataOut[2550]),
.io_dataOut_2551(dataOut[2551]),
.io_dataOut_2552(dataOut[2552]),
.io_dataOut_2553(dataOut[2553]),
.io_dataOut_2554(dataOut[2554]),
.io_dataOut_2555(dataOut[2555]),
.io_dataOut_2556(dataOut[2556]),
.io_dataOut_2557(dataOut[2557]),
.io_dataOut_2558(dataOut[2558]),
.io_dataOut_2559(dataOut[2559]),
.io_dataOut_2560(dataOut[2560]),
.io_dataOut_2561(dataOut[2561]),
.io_dataOut_2562(dataOut[2562]),
.io_dataOut_2563(dataOut[2563]),
.io_dataOut_2564(dataOut[2564]),
.io_dataOut_2565(dataOut[2565]),
.io_dataOut_2566(dataOut[2566]),
.io_dataOut_2567(dataOut[2567]),
.io_dataOut_2568(dataOut[2568]),
.io_dataOut_2569(dataOut[2569]),
.io_dataOut_2570(dataOut[2570]),
.io_dataOut_2571(dataOut[2571]),
.io_dataOut_2572(dataOut[2572]),
.io_dataOut_2573(dataOut[2573]),
.io_dataOut_2574(dataOut[2574]),
.io_dataOut_2575(dataOut[2575]),
.io_dataOut_2576(dataOut[2576]),
.io_dataOut_2577(dataOut[2577]),
.io_dataOut_2578(dataOut[2578]),
.io_dataOut_2579(dataOut[2579]),
.io_dataOut_2580(dataOut[2580]),
.io_dataOut_2581(dataOut[2581]),
.io_dataOut_2582(dataOut[2582]),
.io_dataOut_2583(dataOut[2583]),
.io_dataOut_2584(dataOut[2584]),
.io_dataOut_2585(dataOut[2585]),
.io_dataOut_2586(dataOut[2586]),
.io_dataOut_2587(dataOut[2587]),
.io_dataOut_2588(dataOut[2588]),
.io_dataOut_2589(dataOut[2589]),
.io_dataOut_2590(dataOut[2590]),
.io_dataOut_2591(dataOut[2591]),
.io_dataOut_2592(dataOut[2592]),
.io_dataOut_2593(dataOut[2593]),
.io_dataOut_2594(dataOut[2594]),
.io_dataOut_2595(dataOut[2595]),
.io_dataOut_2596(dataOut[2596]),
.io_dataOut_2597(dataOut[2597]),
.io_dataOut_2598(dataOut[2598]),
.io_dataOut_2599(dataOut[2599]),
.io_dataOut_2600(dataOut[2600]),
.io_dataOut_2601(dataOut[2601]),
.io_dataOut_2602(dataOut[2602]),
.io_dataOut_2603(dataOut[2603]),
.io_dataOut_2604(dataOut[2604]),
.io_dataOut_2605(dataOut[2605]),
.io_dataOut_2606(dataOut[2606]),
.io_dataOut_2607(dataOut[2607]),
.io_dataOut_2608(dataOut[2608]),
.io_dataOut_2609(dataOut[2609]),
.io_dataOut_2610(dataOut[2610]),
.io_dataOut_2611(dataOut[2611]),
.io_dataOut_2612(dataOut[2612]),
.io_dataOut_2613(dataOut[2613]),
.io_dataOut_2614(dataOut[2614]),
.io_dataOut_2615(dataOut[2615]),
.io_dataOut_2616(dataOut[2616]),
.io_dataOut_2617(dataOut[2617]),
.io_dataOut_2618(dataOut[2618]),
.io_dataOut_2619(dataOut[2619]),
.io_dataOut_2620(dataOut[2620]),
.io_dataOut_2621(dataOut[2621]),
.io_dataOut_2622(dataOut[2622]),
.io_dataOut_2623(dataOut[2623]),
.io_dataOut_2624(dataOut[2624]),
.io_dataOut_2625(dataOut[2625]),
.io_dataOut_2626(dataOut[2626]),
.io_dataOut_2627(dataOut[2627]),
.io_dataOut_2628(dataOut[2628]),
.io_dataOut_2629(dataOut[2629]),
.io_dataOut_2630(dataOut[2630]),
.io_dataOut_2631(dataOut[2631]),
.io_dataOut_2632(dataOut[2632]),
.io_dataOut_2633(dataOut[2633]),
.io_dataOut_2634(dataOut[2634]),
.io_dataOut_2635(dataOut[2635]),
.io_dataOut_2636(dataOut[2636]),
.io_dataOut_2637(dataOut[2637]),
.io_dataOut_2638(dataOut[2638]),
.io_dataOut_2639(dataOut[2639]),
.io_dataOut_2640(dataOut[2640]),
.io_dataOut_2641(dataOut[2641]),
.io_dataOut_2642(dataOut[2642]),
.io_dataOut_2643(dataOut[2643]),
.io_dataOut_2644(dataOut[2644]),
.io_dataOut_2645(dataOut[2645]),
.io_dataOut_2646(dataOut[2646]),
.io_dataOut_2647(dataOut[2647]),
.io_dataOut_2648(dataOut[2648]),
.io_dataOut_2649(dataOut[2649]),
.io_dataOut_2650(dataOut[2650]),
.io_dataOut_2651(dataOut[2651]),
.io_dataOut_2652(dataOut[2652]),
.io_dataOut_2653(dataOut[2653]),
.io_dataOut_2654(dataOut[2654]),
.io_dataOut_2655(dataOut[2655]),
.io_dataOut_2656(dataOut[2656]),
.io_dataOut_2657(dataOut[2657]),
.io_dataOut_2658(dataOut[2658]),
.io_dataOut_2659(dataOut[2659]),
.io_dataOut_2660(dataOut[2660]),
.io_dataOut_2661(dataOut[2661]),
.io_dataOut_2662(dataOut[2662]),
.io_dataOut_2663(dataOut[2663]),
.io_dataOut_2664(dataOut[2664]),
.io_dataOut_2665(dataOut[2665]),
.io_dataOut_2666(dataOut[2666]),
.io_dataOut_2667(dataOut[2667]),
.io_dataOut_2668(dataOut[2668]),
.io_dataOut_2669(dataOut[2669]),
.io_dataOut_2670(dataOut[2670]),
.io_dataOut_2671(dataOut[2671]),
.io_dataOut_2672(dataOut[2672]),
.io_dataOut_2673(dataOut[2673]),
.io_dataOut_2674(dataOut[2674]),
.io_dataOut_2675(dataOut[2675]),
.io_dataOut_2676(dataOut[2676]),
.io_dataOut_2677(dataOut[2677]),
.io_dataOut_2678(dataOut[2678]),
.io_dataOut_2679(dataOut[2679]),
.io_dataOut_2680(dataOut[2680]),
.io_dataOut_2681(dataOut[2681]),
.io_dataOut_2682(dataOut[2682]),
.io_dataOut_2683(dataOut[2683]),
.io_dataOut_2684(dataOut[2684]),
.io_dataOut_2685(dataOut[2685]),
.io_dataOut_2686(dataOut[2686]),
.io_dataOut_2687(dataOut[2687]),
.io_dataOut_2688(dataOut[2688]),
.io_dataOut_2689(dataOut[2689]),
.io_dataOut_2690(dataOut[2690]),
.io_dataOut_2691(dataOut[2691]),
.io_dataOut_2692(dataOut[2692]),
.io_dataOut_2693(dataOut[2693]),
.io_dataOut_2694(dataOut[2694]),
.io_dataOut_2695(dataOut[2695]),
.io_dataOut_2696(dataOut[2696]),
.io_dataOut_2697(dataOut[2697]),
.io_dataOut_2698(dataOut[2698]),
.io_dataOut_2699(dataOut[2699]),
.io_dataOut_2700(dataOut[2700]),
.io_dataOut_2701(dataOut[2701]),
.io_dataOut_2702(dataOut[2702]),
.io_dataOut_2703(dataOut[2703]),
.io_dataOut_2704(dataOut[2704]),
.io_dataOut_2705(dataOut[2705]),
.io_dataOut_2706(dataOut[2706]),
.io_dataOut_2707(dataOut[2707]),
.io_dataOut_2708(dataOut[2708]),
.io_dataOut_2709(dataOut[2709]),
.io_dataOut_2710(dataOut[2710]),
.io_dataOut_2711(dataOut[2711]),
.io_dataOut_2712(dataOut[2712]),
.io_dataOut_2713(dataOut[2713]),
.io_dataOut_2714(dataOut[2714]),
.io_dataOut_2715(dataOut[2715]),
.io_dataOut_2716(dataOut[2716]),
.io_dataOut_2717(dataOut[2717]),
.io_dataOut_2718(dataOut[2718]),
.io_dataOut_2719(dataOut[2719]),
.io_dataOut_2720(dataOut[2720]),
.io_dataOut_2721(dataOut[2721]),
.io_dataOut_2722(dataOut[2722]),
.io_dataOut_2723(dataOut[2723]),
.io_dataOut_2724(dataOut[2724]),
.io_dataOut_2725(dataOut[2725]),
.io_dataOut_2726(dataOut[2726]),
.io_dataOut_2727(dataOut[2727]),
.io_dataOut_2728(dataOut[2728]),
.io_dataOut_2729(dataOut[2729]),
.io_dataOut_2730(dataOut[2730]),
.io_dataOut_2731(dataOut[2731]),
.io_dataOut_2732(dataOut[2732]),
.io_dataOut_2733(dataOut[2733]),
.io_dataOut_2734(dataOut[2734]),
.io_dataOut_2735(dataOut[2735]),
.io_dataOut_2736(dataOut[2736]),
.io_dataOut_2737(dataOut[2737]),
.io_dataOut_2738(dataOut[2738]),
.io_dataOut_2739(dataOut[2739]),
.io_dataOut_2740(dataOut[2740]),
.io_dataOut_2741(dataOut[2741]),
.io_dataOut_2742(dataOut[2742]),
.io_dataOut_2743(dataOut[2743]),
.io_dataOut_2744(dataOut[2744]),
.io_dataOut_2745(dataOut[2745]),
.io_dataOut_2746(dataOut[2746]),
.io_dataOut_2747(dataOut[2747]),
.io_dataOut_2748(dataOut[2748]),
.io_dataOut_2749(dataOut[2749]),
.io_dataOut_2750(dataOut[2750]),
.io_dataOut_2751(dataOut[2751]),
.io_dataOut_2752(dataOut[2752]),
.io_dataOut_2753(dataOut[2753]),
.io_dataOut_2754(dataOut[2754]),
.io_dataOut_2755(dataOut[2755]),
.io_dataOut_2756(dataOut[2756]),
.io_dataOut_2757(dataOut[2757]),
.io_dataOut_2758(dataOut[2758]),
.io_dataOut_2759(dataOut[2759]),
.io_dataOut_2760(dataOut[2760]),
.io_dataOut_2761(dataOut[2761]),
.io_dataOut_2762(dataOut[2762]),
.io_dataOut_2763(dataOut[2763]),
.io_dataOut_2764(dataOut[2764]),
.io_dataOut_2765(dataOut[2765]),
.io_dataOut_2766(dataOut[2766]),
.io_dataOut_2767(dataOut[2767]),
.io_dataOut_2768(dataOut[2768]),
.io_dataOut_2769(dataOut[2769]),
.io_dataOut_2770(dataOut[2770]),
.io_dataOut_2771(dataOut[2771]),
.io_dataOut_2772(dataOut[2772]),
.io_dataOut_2773(dataOut[2773]),
.io_dataOut_2774(dataOut[2774]),
.io_dataOut_2775(dataOut[2775]),
.io_dataOut_2776(dataOut[2776]),
.io_dataOut_2777(dataOut[2777]),
.io_dataOut_2778(dataOut[2778]),
.io_dataOut_2779(dataOut[2779]),
.io_dataOut_2780(dataOut[2780]),
.io_dataOut_2781(dataOut[2781]),
.io_dataOut_2782(dataOut[2782]),
.io_dataOut_2783(dataOut[2783]),
.io_dataOut_2784(dataOut[2784]),
.io_dataOut_2785(dataOut[2785]),
.io_dataOut_2786(dataOut[2786]),
.io_dataOut_2787(dataOut[2787]),
.io_dataOut_2788(dataOut[2788]),
.io_dataOut_2789(dataOut[2789]),
.io_dataOut_2790(dataOut[2790]),
.io_dataOut_2791(dataOut[2791]),
.io_dataOut_2792(dataOut[2792]),
.io_dataOut_2793(dataOut[2793]),
.io_dataOut_2794(dataOut[2794]),
.io_dataOut_2795(dataOut[2795]),
.io_dataOut_2796(dataOut[2796]),
.io_dataOut_2797(dataOut[2797]),
.io_dataOut_2798(dataOut[2798]),
.io_dataOut_2799(dataOut[2799]),
.io_dataOut_2800(dataOut[2800]),
.io_dataOut_2801(dataOut[2801]),
.io_dataOut_2802(dataOut[2802]),
.io_dataOut_2803(dataOut[2803]),
.io_dataOut_2804(dataOut[2804]),
.io_dataOut_2805(dataOut[2805]),
.io_dataOut_2806(dataOut[2806]),
.io_dataOut_2807(dataOut[2807]),
.io_dataOut_2808(dataOut[2808]),
.io_dataOut_2809(dataOut[2809]),
.io_dataOut_2810(dataOut[2810]),
.io_dataOut_2811(dataOut[2811]),
.io_dataOut_2812(dataOut[2812]),
.io_dataOut_2813(dataOut[2813]),
.io_dataOut_2814(dataOut[2814]),
.io_dataOut_2815(dataOut[2815]),
.io_dataOut_2816(dataOut[2816]),
.io_dataOut_2817(dataOut[2817]),
.io_dataOut_2818(dataOut[2818]),
.io_dataOut_2819(dataOut[2819]),
.io_dataOut_2820(dataOut[2820]),
.io_dataOut_2821(dataOut[2821]),
.io_dataOut_2822(dataOut[2822]),
.io_dataOut_2823(dataOut[2823]),
.io_dataOut_2824(dataOut[2824]),
.io_dataOut_2825(dataOut[2825]),
.io_dataOut_2826(dataOut[2826]),
.io_dataOut_2827(dataOut[2827]),
.io_dataOut_2828(dataOut[2828]),
.io_dataOut_2829(dataOut[2829]),
.io_dataOut_2830(dataOut[2830]),
.io_dataOut_2831(dataOut[2831]),
.io_dataOut_2832(dataOut[2832]),
.io_dataOut_2833(dataOut[2833]),
.io_dataOut_2834(dataOut[2834]),
.io_dataOut_2835(dataOut[2835]),
.io_dataOut_2836(dataOut[2836]),
.io_dataOut_2837(dataOut[2837]),
.io_dataOut_2838(dataOut[2838]),
.io_dataOut_2839(dataOut[2839]),
.io_dataOut_2840(dataOut[2840]),
.io_dataOut_2841(dataOut[2841]),
.io_dataOut_2842(dataOut[2842]),
.io_dataOut_2843(dataOut[2843]),
.io_dataOut_2844(dataOut[2844]),
.io_dataOut_2845(dataOut[2845]),
.io_dataOut_2846(dataOut[2846]),
.io_dataOut_2847(dataOut[2847]),
.io_dataOut_2848(dataOut[2848]),
.io_dataOut_2849(dataOut[2849]),
.io_dataOut_2850(dataOut[2850]),
.io_dataOut_2851(dataOut[2851]),
.io_dataOut_2852(dataOut[2852]),
.io_dataOut_2853(dataOut[2853]),
.io_dataOut_2854(dataOut[2854]),
.io_dataOut_2855(dataOut[2855]),
.io_dataOut_2856(dataOut[2856]),
.io_dataOut_2857(dataOut[2857]),
.io_dataOut_2858(dataOut[2858]),
.io_dataOut_2859(dataOut[2859]),
.io_dataOut_2860(dataOut[2860]),
.io_dataOut_2861(dataOut[2861]),
.io_dataOut_2862(dataOut[2862]),
.io_dataOut_2863(dataOut[2863]),
.io_dataOut_2864(dataOut[2864]),
.io_dataOut_2865(dataOut[2865]),
.io_dataOut_2866(dataOut[2866]),
.io_dataOut_2867(dataOut[2867]),
.io_dataOut_2868(dataOut[2868]),
.io_dataOut_2869(dataOut[2869]),
.io_dataOut_2870(dataOut[2870]),
.io_dataOut_2871(dataOut[2871]),
.io_dataOut_2872(dataOut[2872]),
.io_dataOut_2873(dataOut[2873]),
.io_dataOut_2874(dataOut[2874]),
.io_dataOut_2875(dataOut[2875]),
.io_dataOut_2876(dataOut[2876]),
.io_dataOut_2877(dataOut[2877]),
.io_dataOut_2878(dataOut[2878]),
.io_dataOut_2879(dataOut[2879]),
.io_dataOut_2880(dataOut[2880]),
.io_dataOut_2881(dataOut[2881]),
.io_dataOut_2882(dataOut[2882]),
.io_dataOut_2883(dataOut[2883]),
.io_dataOut_2884(dataOut[2884]),
.io_dataOut_2885(dataOut[2885]),
.io_dataOut_2886(dataOut[2886]),
.io_dataOut_2887(dataOut[2887]),
.io_dataOut_2888(dataOut[2888]),
.io_dataOut_2889(dataOut[2889]),
.io_dataOut_2890(dataOut[2890]),
.io_dataOut_2891(dataOut[2891]),
.io_dataOut_2892(dataOut[2892]),
.io_dataOut_2893(dataOut[2893]),
.io_dataOut_2894(dataOut[2894]),
.io_dataOut_2895(dataOut[2895]),
.io_dataOut_2896(dataOut[2896]),
.io_dataOut_2897(dataOut[2897]),
.io_dataOut_2898(dataOut[2898]),
.io_dataOut_2899(dataOut[2899]),
.io_dataOut_2900(dataOut[2900]),
.io_dataOut_2901(dataOut[2901]),
.io_dataOut_2902(dataOut[2902]),
.io_dataOut_2903(dataOut[2903]),
.io_dataOut_2904(dataOut[2904]),
.io_dataOut_2905(dataOut[2905]),
.io_dataOut_2906(dataOut[2906]),
.io_dataOut_2907(dataOut[2907]),
.io_dataOut_2908(dataOut[2908]),
.io_dataOut_2909(dataOut[2909]),
.io_dataOut_2910(dataOut[2910]),
.io_dataOut_2911(dataOut[2911]),
.io_dataOut_2912(dataOut[2912]),
.io_dataOut_2913(dataOut[2913]),
.io_dataOut_2914(dataOut[2914]),
.io_dataOut_2915(dataOut[2915]),
.io_dataOut_2916(dataOut[2916]),
.io_dataOut_2917(dataOut[2917]),
.io_dataOut_2918(dataOut[2918]),
.io_dataOut_2919(dataOut[2919]),
.io_dataOut_2920(dataOut[2920]),
.io_dataOut_2921(dataOut[2921]),
.io_dataOut_2922(dataOut[2922]),
.io_dataOut_2923(dataOut[2923]),
.io_dataOut_2924(dataOut[2924]),
.io_dataOut_2925(dataOut[2925]),
.io_dataOut_2926(dataOut[2926]),
.io_dataOut_2927(dataOut[2927]),
.io_dataOut_2928(dataOut[2928]),
.io_dataOut_2929(dataOut[2929]),
.io_dataOut_2930(dataOut[2930]),
.io_dataOut_2931(dataOut[2931]),
.io_dataOut_2932(dataOut[2932]),
.io_dataOut_2933(dataOut[2933]),
.io_dataOut_2934(dataOut[2934]),
.io_dataOut_2935(dataOut[2935]),
.io_dataOut_2936(dataOut[2936]),
.io_dataOut_2937(dataOut[2937]),
.io_dataOut_2938(dataOut[2938]),
.io_dataOut_2939(dataOut[2939]),
.io_dataOut_2940(dataOut[2940]),
.io_dataOut_2941(dataOut[2941]),
.io_dataOut_2942(dataOut[2942]),
.io_dataOut_2943(dataOut[2943]),
.io_dataOut_2944(dataOut[2944]),
.io_dataOut_2945(dataOut[2945]),
.io_dataOut_2946(dataOut[2946]),
.io_dataOut_2947(dataOut[2947]),
.io_dataOut_2948(dataOut[2948]),
.io_dataOut_2949(dataOut[2949]),
.io_dataOut_2950(dataOut[2950]),
.io_dataOut_2951(dataOut[2951]),
.io_dataOut_2952(dataOut[2952]),
.io_dataOut_2953(dataOut[2953]),
.io_dataOut_2954(dataOut[2954]),
.io_dataOut_2955(dataOut[2955]),
.io_dataOut_2956(dataOut[2956]),
.io_dataOut_2957(dataOut[2957]),
.io_dataOut_2958(dataOut[2958]),
.io_dataOut_2959(dataOut[2959]),
.io_dataOut_2960(dataOut[2960]),
.io_dataOut_2961(dataOut[2961]),
.io_dataOut_2962(dataOut[2962]),
.io_dataOut_2963(dataOut[2963]),
.io_dataOut_2964(dataOut[2964]),
.io_dataOut_2965(dataOut[2965]),
.io_dataOut_2966(dataOut[2966]),
.io_dataOut_2967(dataOut[2967]),
.io_dataOut_2968(dataOut[2968]),
.io_dataOut_2969(dataOut[2969]),
.io_dataOut_2970(dataOut[2970]),
.io_dataOut_2971(dataOut[2971]),
.io_dataOut_2972(dataOut[2972]),
.io_dataOut_2973(dataOut[2973]),
.io_dataOut_2974(dataOut[2974]),
.io_dataOut_2975(dataOut[2975]),
.io_dataOut_2976(dataOut[2976]),
.io_dataOut_2977(dataOut[2977]),
.io_dataOut_2978(dataOut[2978]),
.io_dataOut_2979(dataOut[2979]),
.io_dataOut_2980(dataOut[2980]),
.io_dataOut_2981(dataOut[2981]),
.io_dataOut_2982(dataOut[2982]),
.io_dataOut_2983(dataOut[2983]),
.io_dataOut_2984(dataOut[2984]),
.io_dataOut_2985(dataOut[2985]),
.io_dataOut_2986(dataOut[2986]),
.io_dataOut_2987(dataOut[2987]),
.io_dataOut_2988(dataOut[2988]),
.io_dataOut_2989(dataOut[2989]),
.io_dataOut_2990(dataOut[2990]),
.io_dataOut_2991(dataOut[2991]),
.io_dataOut_2992(dataOut[2992]),
.io_dataOut_2993(dataOut[2993]),
.io_dataOut_2994(dataOut[2994]),
.io_dataOut_2995(dataOut[2995]),
.io_dataOut_2996(dataOut[2996]),
.io_dataOut_2997(dataOut[2997]),
.io_dataOut_2998(dataOut[2998]),
.io_dataOut_2999(dataOut[2999]),
.io_dataOut_3000(dataOut[3000]),
.io_dataOut_3001(dataOut[3001]),
.io_dataOut_3002(dataOut[3002]),
.io_dataOut_3003(dataOut[3003]),
.io_dataOut_3004(dataOut[3004]),
.io_dataOut_3005(dataOut[3005]),
.io_dataOut_3006(dataOut[3006]),
.io_dataOut_3007(dataOut[3007]),
.io_dataOut_3008(dataOut[3008]),
.io_dataOut_3009(dataOut[3009]),
.io_dataOut_3010(dataOut[3010]),
.io_dataOut_3011(dataOut[3011]),
.io_dataOut_3012(dataOut[3012]),
.io_dataOut_3013(dataOut[3013]),
.io_dataOut_3014(dataOut[3014]),
.io_dataOut_3015(dataOut[3015]),
.io_dataOut_3016(dataOut[3016]),
.io_dataOut_3017(dataOut[3017]),
.io_dataOut_3018(dataOut[3018]),
.io_dataOut_3019(dataOut[3019]),
.io_dataOut_3020(dataOut[3020]),
.io_dataOut_3021(dataOut[3021]),
.io_dataOut_3022(dataOut[3022]),
.io_dataOut_3023(dataOut[3023]),
.io_dataOut_3024(dataOut[3024]),
.io_dataOut_3025(dataOut[3025]),
.io_dataOut_3026(dataOut[3026]),
.io_dataOut_3027(dataOut[3027]),
.io_dataOut_3028(dataOut[3028]),
.io_dataOut_3029(dataOut[3029]),
.io_dataOut_3030(dataOut[3030]),
.io_dataOut_3031(dataOut[3031]),
.io_dataOut_3032(dataOut[3032]),
.io_dataOut_3033(dataOut[3033]),
.io_dataOut_3034(dataOut[3034]),
.io_dataOut_3035(dataOut[3035]),
.io_dataOut_3036(dataOut[3036]),
.io_dataOut_3037(dataOut[3037]),
.io_dataOut_3038(dataOut[3038]),
.io_dataOut_3039(dataOut[3039]),
.io_dataOut_3040(dataOut[3040]),
.io_dataOut_3041(dataOut[3041]),
.io_dataOut_3042(dataOut[3042]),
.io_dataOut_3043(dataOut[3043]),
.io_dataOut_3044(dataOut[3044]),
.io_dataOut_3045(dataOut[3045]),
.io_dataOut_3046(dataOut[3046]),
.io_dataOut_3047(dataOut[3047]),
.io_dataOut_3048(dataOut[3048]),
.io_dataOut_3049(dataOut[3049]),
.io_dataOut_3050(dataOut[3050]),
.io_dataOut_3051(dataOut[3051]),
.io_dataOut_3052(dataOut[3052]),
.io_dataOut_3053(dataOut[3053]),
.io_dataOut_3054(dataOut[3054]),
.io_dataOut_3055(dataOut[3055]),
.io_dataOut_3056(dataOut[3056]),
.io_dataOut_3057(dataOut[3057]),
.io_dataOut_3058(dataOut[3058]),
.io_dataOut_3059(dataOut[3059]),
.io_dataOut_3060(dataOut[3060]),
.io_dataOut_3061(dataOut[3061]),
.io_dataOut_3062(dataOut[3062]),
.io_dataOut_3063(dataOut[3063]),
.io_dataOut_3064(dataOut[3064]),
.io_dataOut_3065(dataOut[3065]),
.io_dataOut_3066(dataOut[3066]),
.io_dataOut_3067(dataOut[3067]),
.io_dataOut_3068(dataOut[3068]),
.io_dataOut_3069(dataOut[3069]),
.io_dataOut_3070(dataOut[3070]),
.io_dataOut_3071(dataOut[3071]),
.io_dataOut_3072(dataOut[3072]),
.io_dataOut_3073(dataOut[3073]),
.io_dataOut_3074(dataOut[3074]),
.io_dataOut_3075(dataOut[3075]),
.io_dataOut_3076(dataOut[3076]),
.io_dataOut_3077(dataOut[3077]),
.io_dataOut_3078(dataOut[3078]),
.io_dataOut_3079(dataOut[3079]),
.io_dataOut_3080(dataOut[3080]),
.io_dataOut_3081(dataOut[3081]),
.io_dataOut_3082(dataOut[3082]),
.io_dataOut_3083(dataOut[3083]),
.io_dataOut_3084(dataOut[3084]),
.io_dataOut_3085(dataOut[3085]),
.io_dataOut_3086(dataOut[3086]),
.io_dataOut_3087(dataOut[3087]),
.io_dataOut_3088(dataOut[3088]),
.io_dataOut_3089(dataOut[3089]),
.io_dataOut_3090(dataOut[3090]),
.io_dataOut_3091(dataOut[3091]),
.io_dataOut_3092(dataOut[3092]),
.io_dataOut_3093(dataOut[3093]),
.io_dataOut_3094(dataOut[3094]),
.io_dataOut_3095(dataOut[3095]),
.io_dataOut_3096(dataOut[3096]),
.io_dataOut_3097(dataOut[3097]),
.io_dataOut_3098(dataOut[3098]),
.io_dataOut_3099(dataOut[3099]),
.io_dataOut_3100(dataOut[3100]),
.io_dataOut_3101(dataOut[3101]),
.io_dataOut_3102(dataOut[3102]),
.io_dataOut_3103(dataOut[3103]),
.io_dataOut_3104(dataOut[3104]),
.io_dataOut_3105(dataOut[3105]),
.io_dataOut_3106(dataOut[3106]),
.io_dataOut_3107(dataOut[3107]),
.io_dataOut_3108(dataOut[3108]),
.io_dataOut_3109(dataOut[3109]),
.io_dataOut_3110(dataOut[3110]),
.io_dataOut_3111(dataOut[3111]),
.io_dataOut_3112(dataOut[3112]),
.io_dataOut_3113(dataOut[3113]),
.io_dataOut_3114(dataOut[3114]),
.io_dataOut_3115(dataOut[3115]),
.io_dataOut_3116(dataOut[3116]),
.io_dataOut_3117(dataOut[3117]),
.io_dataOut_3118(dataOut[3118]),
.io_dataOut_3119(dataOut[3119]),
.io_dataOut_3120(dataOut[3120]),
.io_dataOut_3121(dataOut[3121]),
.io_dataOut_3122(dataOut[3122]),
.io_dataOut_3123(dataOut[3123]),
.io_dataOut_3124(dataOut[3124]),
.io_dataOut_3125(dataOut[3125]),
.io_dataOut_3126(dataOut[3126]),
.io_dataOut_3127(dataOut[3127]),
.io_dataOut_3128(dataOut[3128]),
.io_dataOut_3129(dataOut[3129]),
.io_dataOut_3130(dataOut[3130]),
.io_dataOut_3131(dataOut[3131]),
.io_dataOut_3132(dataOut[3132]),
.io_dataOut_3133(dataOut[3133]),
.io_dataOut_3134(dataOut[3134]),
.io_dataOut_3135(dataOut[3135]),
.io_dataOut_3136(dataOut[3136]),
.io_dataOut_3137(dataOut[3137]),
.io_dataOut_3138(dataOut[3138]),
.io_dataOut_3139(dataOut[3139]),
.io_dataOut_3140(dataOut[3140]),
.io_dataOut_3141(dataOut[3141]),
.io_dataOut_3142(dataOut[3142]),
.io_dataOut_3143(dataOut[3143]),
.io_dataOut_3144(dataOut[3144]),
.io_dataOut_3145(dataOut[3145]),
.io_dataOut_3146(dataOut[3146]),
.io_dataOut_3147(dataOut[3147]),
.io_dataOut_3148(dataOut[3148]),
.io_dataOut_3149(dataOut[3149]),
.io_dataOut_3150(dataOut[3150]),
.io_dataOut_3151(dataOut[3151]),
.io_dataOut_3152(dataOut[3152]),
.io_dataOut_3153(dataOut[3153]),
.io_dataOut_3154(dataOut[3154]),
.io_dataOut_3155(dataOut[3155]),
.io_dataOut_3156(dataOut[3156]),
.io_dataOut_3157(dataOut[3157]),
.io_dataOut_3158(dataOut[3158]),
.io_dataOut_3159(dataOut[3159]),
.io_dataOut_3160(dataOut[3160]),
.io_dataOut_3161(dataOut[3161]),
.io_dataOut_3162(dataOut[3162]),
.io_dataOut_3163(dataOut[3163]),
.io_dataOut_3164(dataOut[3164]),
.io_dataOut_3165(dataOut[3165]),
.io_dataOut_3166(dataOut[3166]),
.io_dataOut_3167(dataOut[3167]),
.io_dataOut_3168(dataOut[3168]),
.io_dataOut_3169(dataOut[3169]),
.io_dataOut_3170(dataOut[3170]),
.io_dataOut_3171(dataOut[3171]),
.io_dataOut_3172(dataOut[3172]),
.io_dataOut_3173(dataOut[3173]),
.io_dataOut_3174(dataOut[3174]),
.io_dataOut_3175(dataOut[3175]),
.io_dataOut_3176(dataOut[3176]),
.io_dataOut_3177(dataOut[3177]),
.io_dataOut_3178(dataOut[3178]),
.io_dataOut_3179(dataOut[3179]),
.io_dataOut_3180(dataOut[3180]),
.io_dataOut_3181(dataOut[3181]),
.io_dataOut_3182(dataOut[3182]),
.io_dataOut_3183(dataOut[3183]),
.io_dataOut_3184(dataOut[3184]),
.io_dataOut_3185(dataOut[3185]),
.io_dataOut_3186(dataOut[3186]),
.io_dataOut_3187(dataOut[3187]),
.io_dataOut_3188(dataOut[3188]),
.io_dataOut_3189(dataOut[3189]),
.io_dataOut_3190(dataOut[3190]),
.io_dataOut_3191(dataOut[3191]),
.io_dataOut_3192(dataOut[3192]),
.io_dataOut_3193(dataOut[3193]),
.io_dataOut_3194(dataOut[3194]),
.io_dataOut_3195(dataOut[3195]),
.io_dataOut_3196(dataOut[3196]),
.io_dataOut_3197(dataOut[3197]),
.io_dataOut_3198(dataOut[3198]),
.io_dataOut_3199(dataOut[3199]),
.io_dataOut_3200(dataOut[3200]),
.io_dataOut_3201(dataOut[3201]),
.io_dataOut_3202(dataOut[3202]),
.io_dataOut_3203(dataOut[3203]),
.io_dataOut_3204(dataOut[3204]),
.io_dataOut_3205(dataOut[3205]),
.io_dataOut_3206(dataOut[3206]),
.io_dataOut_3207(dataOut[3207]),
.io_dataOut_3208(dataOut[3208]),
.io_dataOut_3209(dataOut[3209]),
.io_dataOut_3210(dataOut[3210]),
.io_dataOut_3211(dataOut[3211]),
.io_dataOut_3212(dataOut[3212]),
.io_dataOut_3213(dataOut[3213]),
.io_dataOut_3214(dataOut[3214]),
.io_dataOut_3215(dataOut[3215]),
.io_dataOut_3216(dataOut[3216]),
.io_dataOut_3217(dataOut[3217]),
.io_dataOut_3218(dataOut[3218]),
.io_dataOut_3219(dataOut[3219]),
.io_dataOut_3220(dataOut[3220]),
.io_dataOut_3221(dataOut[3221]),
.io_dataOut_3222(dataOut[3222]),
.io_dataOut_3223(dataOut[3223]),
.io_dataOut_3224(dataOut[3224]),
.io_dataOut_3225(dataOut[3225]),
.io_dataOut_3226(dataOut[3226]),
.io_dataOut_3227(dataOut[3227]),
.io_dataOut_3228(dataOut[3228]),
.io_dataOut_3229(dataOut[3229]),
.io_dataOut_3230(dataOut[3230]),
.io_dataOut_3231(dataOut[3231]),
.io_dataOut_3232(dataOut[3232]),
.io_dataOut_3233(dataOut[3233]),
.io_dataOut_3234(dataOut[3234]),
.io_dataOut_3235(dataOut[3235]),
.io_dataOut_3236(dataOut[3236]),
.io_dataOut_3237(dataOut[3237]),
.io_dataOut_3238(dataOut[3238]),
.io_dataOut_3239(dataOut[3239]),
.io_dataOut_3240(dataOut[3240]),
.io_dataOut_3241(dataOut[3241]),
.io_dataOut_3242(dataOut[3242]),
.io_dataOut_3243(dataOut[3243]),
.io_dataOut_3244(dataOut[3244]),
.io_dataOut_3245(dataOut[3245]),
.io_dataOut_3246(dataOut[3246]),
.io_dataOut_3247(dataOut[3247]),
.io_dataOut_3248(dataOut[3248]),
.io_dataOut_3249(dataOut[3249]),
.io_dataOut_3250(dataOut[3250]),
.io_dataOut_3251(dataOut[3251]),
.io_dataOut_3252(dataOut[3252]),
.io_dataOut_3253(dataOut[3253]),
.io_dataOut_3254(dataOut[3254]),
.io_dataOut_3255(dataOut[3255]),
.io_dataOut_3256(dataOut[3256]),
.io_dataOut_3257(dataOut[3257]),
.io_dataOut_3258(dataOut[3258]),
.io_dataOut_3259(dataOut[3259]),
.io_dataOut_3260(dataOut[3260]),
.io_dataOut_3261(dataOut[3261]),
.io_dataOut_3262(dataOut[3262]),
.io_dataOut_3263(dataOut[3263]),
.io_dataOut_3264(dataOut[3264]),
.io_dataOut_3265(dataOut[3265]),
.io_dataOut_3266(dataOut[3266]),
.io_dataOut_3267(dataOut[3267]),
.io_dataOut_3268(dataOut[3268]),
.io_dataOut_3269(dataOut[3269]),
.io_dataOut_3270(dataOut[3270]),
.io_dataOut_3271(dataOut[3271]),
.io_dataOut_3272(dataOut[3272]),
.io_dataOut_3273(dataOut[3273]),
.io_dataOut_3274(dataOut[3274]),
.io_dataOut_3275(dataOut[3275]),
.io_dataOut_3276(dataOut[3276]),
.io_dataOut_3277(dataOut[3277]),
.io_dataOut_3278(dataOut[3278]),
.io_dataOut_3279(dataOut[3279]),
.io_dataOut_3280(dataOut[3280]),
.io_dataOut_3281(dataOut[3281]),
.io_dataOut_3282(dataOut[3282]),
.io_dataOut_3283(dataOut[3283]),
.io_dataOut_3284(dataOut[3284]),
.io_dataOut_3285(dataOut[3285]),
.io_dataOut_3286(dataOut[3286]),
.io_dataOut_3287(dataOut[3287]),
.io_dataOut_3288(dataOut[3288]),
.io_dataOut_3289(dataOut[3289]),
.io_dataOut_3290(dataOut[3290]),
.io_dataOut_3291(dataOut[3291]),
.io_dataOut_3292(dataOut[3292]),
.io_dataOut_3293(dataOut[3293]),
.io_dataOut_3294(dataOut[3294]),
.io_dataOut_3295(dataOut[3295]),
.io_dataOut_3296(dataOut[3296]),
.io_dataOut_3297(dataOut[3297]),
.io_dataOut_3298(dataOut[3298]),
.io_dataOut_3299(dataOut[3299]),
.io_dataOut_3300(dataOut[3300]),
.io_dataOut_3301(dataOut[3301]),
.io_dataOut_3302(dataOut[3302]),
.io_dataOut_3303(dataOut[3303]),
.io_dataOut_3304(dataOut[3304]),
.io_dataOut_3305(dataOut[3305]),
.io_dataOut_3306(dataOut[3306]),
.io_dataOut_3307(dataOut[3307]),
.io_dataOut_3308(dataOut[3308]),
.io_dataOut_3309(dataOut[3309]),
.io_dataOut_3310(dataOut[3310]),
.io_dataOut_3311(dataOut[3311]),
.io_dataOut_3312(dataOut[3312]),
.io_dataOut_3313(dataOut[3313]),
.io_dataOut_3314(dataOut[3314]),
.io_dataOut_3315(dataOut[3315]),
.io_dataOut_3316(dataOut[3316]),
.io_dataOut_3317(dataOut[3317]),
.io_dataOut_3318(dataOut[3318]),
.io_dataOut_3319(dataOut[3319]),
.io_dataOut_3320(dataOut[3320]),
.io_dataOut_3321(dataOut[3321]),
.io_dataOut_3322(dataOut[3322]),
.io_dataOut_3323(dataOut[3323]),
.io_dataOut_3324(dataOut[3324]),
.io_dataOut_3325(dataOut[3325]),
.io_dataOut_3326(dataOut[3326]),
.io_dataOut_3327(dataOut[3327]),
.io_dataOut_3328(dataOut[3328]),
.io_dataOut_3329(dataOut[3329]),
.io_dataOut_3330(dataOut[3330]),
.io_dataOut_3331(dataOut[3331]),
.io_dataOut_3332(dataOut[3332]),
.io_dataOut_3333(dataOut[3333]),
.io_dataOut_3334(dataOut[3334]),
.io_dataOut_3335(dataOut[3335]),
.io_dataOut_3336(dataOut[3336]),
.io_dataOut_3337(dataOut[3337]),
.io_dataOut_3338(dataOut[3338]),
.io_dataOut_3339(dataOut[3339]),
.io_dataOut_3340(dataOut[3340]),
.io_dataOut_3341(dataOut[3341]),
.io_dataOut_3342(dataOut[3342]),
.io_dataOut_3343(dataOut[3343]),
.io_dataOut_3344(dataOut[3344]),
.io_dataOut_3345(dataOut[3345]),
.io_dataOut_3346(dataOut[3346]),
.io_dataOut_3347(dataOut[3347]),
.io_dataOut_3348(dataOut[3348]),
.io_dataOut_3349(dataOut[3349]),
.io_dataOut_3350(dataOut[3350]),
.io_dataOut_3351(dataOut[3351]),
.io_dataOut_3352(dataOut[3352]),
.io_dataOut_3353(dataOut[3353]),
.io_dataOut_3354(dataOut[3354]),
.io_dataOut_3355(dataOut[3355]),
.io_dataOut_3356(dataOut[3356]),
.io_dataOut_3357(dataOut[3357]),
.io_dataOut_3358(dataOut[3358]),
.io_dataOut_3359(dataOut[3359]),
.io_dataOut_3360(dataOut[3360]),
.io_dataOut_3361(dataOut[3361]),
.io_dataOut_3362(dataOut[3362]),
.io_dataOut_3363(dataOut[3363]),
.io_dataOut_3364(dataOut[3364]),
.io_dataOut_3365(dataOut[3365]),
.io_dataOut_3366(dataOut[3366]),
.io_dataOut_3367(dataOut[3367]),
.io_dataOut_3368(dataOut[3368]),
.io_dataOut_3369(dataOut[3369]),
.io_dataOut_3370(dataOut[3370]),
.io_dataOut_3371(dataOut[3371]),
.io_dataOut_3372(dataOut[3372]),
.io_dataOut_3373(dataOut[3373]),
.io_dataOut_3374(dataOut[3374]),
.io_dataOut_3375(dataOut[3375]),
.io_dataOut_3376(dataOut[3376]),
.io_dataOut_3377(dataOut[3377]),
.io_dataOut_3378(dataOut[3378]),
.io_dataOut_3379(dataOut[3379]),
.io_dataOut_3380(dataOut[3380]),
.io_dataOut_3381(dataOut[3381]),
.io_dataOut_3382(dataOut[3382]),
.io_dataOut_3383(dataOut[3383]),
.io_dataOut_3384(dataOut[3384]),
.io_dataOut_3385(dataOut[3385]),
.io_dataOut_3386(dataOut[3386]),
.io_dataOut_3387(dataOut[3387]),
.io_dataOut_3388(dataOut[3388]),
.io_dataOut_3389(dataOut[3389]),
.io_dataOut_3390(dataOut[3390]),
.io_dataOut_3391(dataOut[3391]),
.io_dataOut_3392(dataOut[3392]),
.io_dataOut_3393(dataOut[3393]),
.io_dataOut_3394(dataOut[3394]),
.io_dataOut_3395(dataOut[3395]),
.io_dataOut_3396(dataOut[3396]),
.io_dataOut_3397(dataOut[3397]),
.io_dataOut_3398(dataOut[3398]),
.io_dataOut_3399(dataOut[3399]),
.io_dataOut_3400(dataOut[3400]),
.io_dataOut_3401(dataOut[3401]),
.io_dataOut_3402(dataOut[3402]),
.io_dataOut_3403(dataOut[3403]),
.io_dataOut_3404(dataOut[3404]),
.io_dataOut_3405(dataOut[3405]),
.io_dataOut_3406(dataOut[3406]),
.io_dataOut_3407(dataOut[3407]),
.io_dataOut_3408(dataOut[3408]),
.io_dataOut_3409(dataOut[3409]),
.io_dataOut_3410(dataOut[3410]),
.io_dataOut_3411(dataOut[3411]),
.io_dataOut_3412(dataOut[3412]),
.io_dataOut_3413(dataOut[3413]),
.io_dataOut_3414(dataOut[3414]),
.io_dataOut_3415(dataOut[3415]),
.io_dataOut_3416(dataOut[3416]),
.io_dataOut_3417(dataOut[3417]),
.io_dataOut_3418(dataOut[3418]),
.io_dataOut_3419(dataOut[3419]),
.io_dataOut_3420(dataOut[3420]),
.io_dataOut_3421(dataOut[3421]),
.io_dataOut_3422(dataOut[3422]),
.io_dataOut_3423(dataOut[3423]),
.io_dataOut_3424(dataOut[3424]),
.io_dataOut_3425(dataOut[3425]),
.io_dataOut_3426(dataOut[3426]),
.io_dataOut_3427(dataOut[3427]),
.io_dataOut_3428(dataOut[3428]),
.io_dataOut_3429(dataOut[3429]),
.io_dataOut_3430(dataOut[3430]),
.io_dataOut_3431(dataOut[3431]),
.io_dataOut_3432(dataOut[3432]),
.io_dataOut_3433(dataOut[3433]),
.io_dataOut_3434(dataOut[3434]),
.io_dataOut_3435(dataOut[3435]),
.io_dataOut_3436(dataOut[3436]),
.io_dataOut_3437(dataOut[3437]),
.io_dataOut_3438(dataOut[3438]),
.io_dataOut_3439(dataOut[3439]),
.io_dataOut_3440(dataOut[3440]),
.io_dataOut_3441(dataOut[3441]),
.io_dataOut_3442(dataOut[3442]),
.io_dataOut_3443(dataOut[3443]),
.io_dataOut_3444(dataOut[3444]),
.io_dataOut_3445(dataOut[3445]),
.io_dataOut_3446(dataOut[3446]),
.io_dataOut_3447(dataOut[3447]),
.io_dataOut_3448(dataOut[3448]),
.io_dataOut_3449(dataOut[3449]),
.io_dataOut_3450(dataOut[3450]),
.io_dataOut_3451(dataOut[3451]),
.io_dataOut_3452(dataOut[3452]),
.io_dataOut_3453(dataOut[3453]),
.io_dataOut_3454(dataOut[3454]),
.io_dataOut_3455(dataOut[3455]),
.io_dataOut_3456(dataOut[3456]),
.io_dataOut_3457(dataOut[3457]),
.io_dataOut_3458(dataOut[3458]),
.io_dataOut_3459(dataOut[3459]),
.io_dataOut_3460(dataOut[3460]),
.io_dataOut_3461(dataOut[3461]),
.io_dataOut_3462(dataOut[3462]),
.io_dataOut_3463(dataOut[3463]),
.io_dataOut_3464(dataOut[3464]),
.io_dataOut_3465(dataOut[3465]),
.io_dataOut_3466(dataOut[3466]),
.io_dataOut_3467(dataOut[3467]),
.io_dataOut_3468(dataOut[3468]),
.io_dataOut_3469(dataOut[3469]),
.io_dataOut_3470(dataOut[3470]),
.io_dataOut_3471(dataOut[3471]),
.io_dataOut_3472(dataOut[3472]),
.io_dataOut_3473(dataOut[3473]),
.io_dataOut_3474(dataOut[3474]),
.io_dataOut_3475(dataOut[3475]),
.io_dataOut_3476(dataOut[3476]),
.io_dataOut_3477(dataOut[3477]),
.io_dataOut_3478(dataOut[3478]),
.io_dataOut_3479(dataOut[3479]),
.io_dataOut_3480(dataOut[3480]),
.io_dataOut_3481(dataOut[3481]),
.io_dataOut_3482(dataOut[3482]),
.io_dataOut_3483(dataOut[3483]),
.io_dataOut_3484(dataOut[3484]),
.io_dataOut_3485(dataOut[3485]),
.io_dataOut_3486(dataOut[3486]),
.io_dataOut_3487(dataOut[3487]),
.io_dataOut_3488(dataOut[3488]),
.io_dataOut_3489(dataOut[3489]),
.io_dataOut_3490(dataOut[3490]),
.io_dataOut_3491(dataOut[3491]),
.io_dataOut_3492(dataOut[3492]),
.io_dataOut_3493(dataOut[3493]),
.io_dataOut_3494(dataOut[3494]),
.io_dataOut_3495(dataOut[3495]),
.io_dataOut_3496(dataOut[3496]),
.io_dataOut_3497(dataOut[3497]),
.io_dataOut_3498(dataOut[3498]),
.io_dataOut_3499(dataOut[3499]),
.io_dataOut_3500(dataOut[3500]),
.io_dataOut_3501(dataOut[3501]),
.io_dataOut_3502(dataOut[3502]),
.io_dataOut_3503(dataOut[3503]),
.io_dataOut_3504(dataOut[3504]),
.io_dataOut_3505(dataOut[3505]),
.io_dataOut_3506(dataOut[3506]),
.io_dataOut_3507(dataOut[3507]),
.io_dataOut_3508(dataOut[3508]),
.io_dataOut_3509(dataOut[3509]),
.io_dataOut_3510(dataOut[3510]),
.io_dataOut_3511(dataOut[3511]),
.io_dataOut_3512(dataOut[3512]),
.io_dataOut_3513(dataOut[3513]),
.io_dataOut_3514(dataOut[3514]),
.io_dataOut_3515(dataOut[3515]),
.io_dataOut_3516(dataOut[3516]),
.io_dataOut_3517(dataOut[3517]),
.io_dataOut_3518(dataOut[3518]),
.io_dataOut_3519(dataOut[3519]),
.io_dataOut_3520(dataOut[3520]),
.io_dataOut_3521(dataOut[3521]),
.io_dataOut_3522(dataOut[3522]),
.io_dataOut_3523(dataOut[3523]),
.io_dataOut_3524(dataOut[3524]),
.io_dataOut_3525(dataOut[3525]),
.io_dataOut_3526(dataOut[3526]),
.io_dataOut_3527(dataOut[3527]),
.io_dataOut_3528(dataOut[3528]),
.io_dataOut_3529(dataOut[3529]),
.io_dataOut_3530(dataOut[3530]),
.io_dataOut_3531(dataOut[3531]),
.io_dataOut_3532(dataOut[3532]),
.io_dataOut_3533(dataOut[3533]),
.io_dataOut_3534(dataOut[3534]),
.io_dataOut_3535(dataOut[3535]),
.io_dataOut_3536(dataOut[3536]),
.io_dataOut_3537(dataOut[3537]),
.io_dataOut_3538(dataOut[3538]),
.io_dataOut_3539(dataOut[3539]),
.io_dataOut_3540(dataOut[3540]),
.io_dataOut_3541(dataOut[3541]),
.io_dataOut_3542(dataOut[3542]),
.io_dataOut_3543(dataOut[3543]),
.io_dataOut_3544(dataOut[3544]),
.io_dataOut_3545(dataOut[3545]),
.io_dataOut_3546(dataOut[3546]),
.io_dataOut_3547(dataOut[3547]),
.io_dataOut_3548(dataOut[3548]),
.io_dataOut_3549(dataOut[3549]),
.io_dataOut_3550(dataOut[3550]),
.io_dataOut_3551(dataOut[3551]),
.io_dataOut_3552(dataOut[3552]),
.io_dataOut_3553(dataOut[3553]),
.io_dataOut_3554(dataOut[3554]),
.io_dataOut_3555(dataOut[3555]),
.io_dataOut_3556(dataOut[3556]),
.io_dataOut_3557(dataOut[3557]),
.io_dataOut_3558(dataOut[3558]),
.io_dataOut_3559(dataOut[3559]),
.io_dataOut_3560(dataOut[3560]),
.io_dataOut_3561(dataOut[3561]),
.io_dataOut_3562(dataOut[3562]),
.io_dataOut_3563(dataOut[3563]),
.io_dataOut_3564(dataOut[3564]),
.io_dataOut_3565(dataOut[3565]),
.io_dataOut_3566(dataOut[3566]),
.io_dataOut_3567(dataOut[3567]),
.io_dataOut_3568(dataOut[3568]),
.io_dataOut_3569(dataOut[3569]),
.io_dataOut_3570(dataOut[3570]),
.io_dataOut_3571(dataOut[3571]),
.io_dataOut_3572(dataOut[3572]),
.io_dataOut_3573(dataOut[3573]),
.io_dataOut_3574(dataOut[3574]),
.io_dataOut_3575(dataOut[3575]),
.io_dataOut_3576(dataOut[3576]),
.io_dataOut_3577(dataOut[3577]),
.io_dataOut_3578(dataOut[3578]),
.io_dataOut_3579(dataOut[3579]),
.io_dataOut_3580(dataOut[3580]),
.io_dataOut_3581(dataOut[3581]),
.io_dataOut_3582(dataOut[3582]),
.io_dataOut_3583(dataOut[3583]),
.io_dataOut_3584(dataOut[3584]),
.io_dataOut_3585(dataOut[3585]),
.io_dataOut_3586(dataOut[3586]),
.io_dataOut_3587(dataOut[3587]),
.io_dataOut_3588(dataOut[3588]),
.io_dataOut_3589(dataOut[3589]),
.io_dataOut_3590(dataOut[3590]),
.io_dataOut_3591(dataOut[3591]),
.io_dataOut_3592(dataOut[3592]),
.io_dataOut_3593(dataOut[3593]),
.io_dataOut_3594(dataOut[3594]),
.io_dataOut_3595(dataOut[3595]),
.io_dataOut_3596(dataOut[3596]),
.io_dataOut_3597(dataOut[3597]),
.io_dataOut_3598(dataOut[3598]),
.io_dataOut_3599(dataOut[3599]),
.io_dataOut_3600(dataOut[3600]),
.io_dataOut_3601(dataOut[3601]),
.io_dataOut_3602(dataOut[3602]),
.io_dataOut_3603(dataOut[3603]),
.io_dataOut_3604(dataOut[3604]),
.io_dataOut_3605(dataOut[3605]),
.io_dataOut_3606(dataOut[3606]),
.io_dataOut_3607(dataOut[3607]),
.io_dataOut_3608(dataOut[3608]),
.io_dataOut_3609(dataOut[3609]),
.io_dataOut_3610(dataOut[3610]),
.io_dataOut_3611(dataOut[3611]),
.io_dataOut_3612(dataOut[3612]),
.io_dataOut_3613(dataOut[3613]),
.io_dataOut_3614(dataOut[3614]),
.io_dataOut_3615(dataOut[3615]),
.io_dataOut_3616(dataOut[3616]),
.io_dataOut_3617(dataOut[3617]),
.io_dataOut_3618(dataOut[3618]),
.io_dataOut_3619(dataOut[3619]),
.io_dataOut_3620(dataOut[3620]),
.io_dataOut_3621(dataOut[3621]),
.io_dataOut_3622(dataOut[3622]),
.io_dataOut_3623(dataOut[3623]),
.io_dataOut_3624(dataOut[3624]),
.io_dataOut_3625(dataOut[3625]),
.io_dataOut_3626(dataOut[3626]),
.io_dataOut_3627(dataOut[3627]),
.io_dataOut_3628(dataOut[3628]),
.io_dataOut_3629(dataOut[3629]),
.io_dataOut_3630(dataOut[3630]),
.io_dataOut_3631(dataOut[3631]),
.io_dataOut_3632(dataOut[3632]),
.io_dataOut_3633(dataOut[3633]),
.io_dataOut_3634(dataOut[3634]),
.io_dataOut_3635(dataOut[3635]),
.io_dataOut_3636(dataOut[3636]),
.io_dataOut_3637(dataOut[3637]),
.io_dataOut_3638(dataOut[3638]),
.io_dataOut_3639(dataOut[3639]),
.io_dataOut_3640(dataOut[3640]),
.io_dataOut_3641(dataOut[3641]),
.io_dataOut_3642(dataOut[3642]),
.io_dataOut_3643(dataOut[3643]),
.io_dataOut_3644(dataOut[3644]),
.io_dataOut_3645(dataOut[3645]),
.io_dataOut_3646(dataOut[3646]),
.io_dataOut_3647(dataOut[3647]),
.io_dataOut_3648(dataOut[3648]),
.io_dataOut_3649(dataOut[3649]),
.io_dataOut_3650(dataOut[3650]),
.io_dataOut_3651(dataOut[3651]),
.io_dataOut_3652(dataOut[3652]),
.io_dataOut_3653(dataOut[3653]),
.io_dataOut_3654(dataOut[3654]),
.io_dataOut_3655(dataOut[3655]),
.io_dataOut_3656(dataOut[3656]),
.io_dataOut_3657(dataOut[3657]),
.io_dataOut_3658(dataOut[3658]),
.io_dataOut_3659(dataOut[3659]),
.io_dataOut_3660(dataOut[3660]),
.io_dataOut_3661(dataOut[3661]),
.io_dataOut_3662(dataOut[3662]),
.io_dataOut_3663(dataOut[3663]),
.io_dataOut_3664(dataOut[3664]),
.io_dataOut_3665(dataOut[3665]),
.io_dataOut_3666(dataOut[3666]),
.io_dataOut_3667(dataOut[3667]),
.io_dataOut_3668(dataOut[3668]),
.io_dataOut_3669(dataOut[3669]),
.io_dataOut_3670(dataOut[3670]),
.io_dataOut_3671(dataOut[3671]),
.io_dataOut_3672(dataOut[3672]),
.io_dataOut_3673(dataOut[3673]),
.io_dataOut_3674(dataOut[3674]),
.io_dataOut_3675(dataOut[3675]),
.io_dataOut_3676(dataOut[3676]),
.io_dataOut_3677(dataOut[3677]),
.io_dataOut_3678(dataOut[3678]),
.io_dataOut_3679(dataOut[3679]),
.io_dataOut_3680(dataOut[3680]),
.io_dataOut_3681(dataOut[3681]),
.io_dataOut_3682(dataOut[3682]),
.io_dataOut_3683(dataOut[3683]),
.io_dataOut_3684(dataOut[3684]),
.io_dataOut_3685(dataOut[3685]),
.io_dataOut_3686(dataOut[3686]),
.io_dataOut_3687(dataOut[3687]),
.io_dataOut_3688(dataOut[3688]),
.io_dataOut_3689(dataOut[3689]),
.io_dataOut_3690(dataOut[3690]),
.io_dataOut_3691(dataOut[3691]),
.io_dataOut_3692(dataOut[3692]),
.io_dataOut_3693(dataOut[3693]),
.io_dataOut_3694(dataOut[3694]),
.io_dataOut_3695(dataOut[3695]),
.io_dataOut_3696(dataOut[3696]),
.io_dataOut_3697(dataOut[3697]),
.io_dataOut_3698(dataOut[3698]),
.io_dataOut_3699(dataOut[3699]),
.io_dataOut_3700(dataOut[3700]),
.io_dataOut_3701(dataOut[3701]),
.io_dataOut_3702(dataOut[3702]),
.io_dataOut_3703(dataOut[3703]),
.io_dataOut_3704(dataOut[3704]),
.io_dataOut_3705(dataOut[3705]),
.io_dataOut_3706(dataOut[3706]),
.io_dataOut_3707(dataOut[3707]),
.io_dataOut_3708(dataOut[3708]),
.io_dataOut_3709(dataOut[3709]),
.io_dataOut_3710(dataOut[3710]),
.io_dataOut_3711(dataOut[3711]),
.io_dataOut_3712(dataOut[3712]),
.io_dataOut_3713(dataOut[3713]),
.io_dataOut_3714(dataOut[3714]),
.io_dataOut_3715(dataOut[3715]),
.io_dataOut_3716(dataOut[3716]),
.io_dataOut_3717(dataOut[3717]),
.io_dataOut_3718(dataOut[3718]),
.io_dataOut_3719(dataOut[3719]),
.io_dataOut_3720(dataOut[3720]),
.io_dataOut_3721(dataOut[3721]),
.io_dataOut_3722(dataOut[3722]),
.io_dataOut_3723(dataOut[3723]),
.io_dataOut_3724(dataOut[3724]),
.io_dataOut_3725(dataOut[3725]),
.io_dataOut_3726(dataOut[3726]),
.io_dataOut_3727(dataOut[3727]),
.io_dataOut_3728(dataOut[3728]),
.io_dataOut_3729(dataOut[3729]),
.io_dataOut_3730(dataOut[3730]),
.io_dataOut_3731(dataOut[3731]),
.io_dataOut_3732(dataOut[3732]),
.io_dataOut_3733(dataOut[3733]),
.io_dataOut_3734(dataOut[3734]),
.io_dataOut_3735(dataOut[3735]),
.io_dataOut_3736(dataOut[3736]),
.io_dataOut_3737(dataOut[3737]),
.io_dataOut_3738(dataOut[3738]),
.io_dataOut_3739(dataOut[3739]),
.io_dataOut_3740(dataOut[3740]),
.io_dataOut_3741(dataOut[3741]),
.io_dataOut_3742(dataOut[3742]),
.io_dataOut_3743(dataOut[3743]),
.io_dataOut_3744(dataOut[3744]),
.io_dataOut_3745(dataOut[3745]),
.io_dataOut_3746(dataOut[3746]),
.io_dataOut_3747(dataOut[3747]),
.io_dataOut_3748(dataOut[3748]),
.io_dataOut_3749(dataOut[3749]),
.io_dataOut_3750(dataOut[3750]),
.io_dataOut_3751(dataOut[3751]),
.io_dataOut_3752(dataOut[3752]),
.io_dataOut_3753(dataOut[3753]),
.io_dataOut_3754(dataOut[3754]),
.io_dataOut_3755(dataOut[3755]),
.io_dataOut_3756(dataOut[3756]),
.io_dataOut_3757(dataOut[3757]),
.io_dataOut_3758(dataOut[3758]),
.io_dataOut_3759(dataOut[3759]),
.io_dataOut_3760(dataOut[3760]),
.io_dataOut_3761(dataOut[3761]),
.io_dataOut_3762(dataOut[3762]),
.io_dataOut_3763(dataOut[3763]),
.io_dataOut_3764(dataOut[3764]),
.io_dataOut_3765(dataOut[3765]),
.io_dataOut_3766(dataOut[3766]),
.io_dataOut_3767(dataOut[3767]),
.io_dataOut_3768(dataOut[3768]),
.io_dataOut_3769(dataOut[3769]),
.io_dataOut_3770(dataOut[3770]),
.io_dataOut_3771(dataOut[3771]),
.io_dataOut_3772(dataOut[3772]),
.io_dataOut_3773(dataOut[3773]),
.io_dataOut_3774(dataOut[3774]),
.io_dataOut_3775(dataOut[3775]),
.io_dataOut_3776(dataOut[3776]),
.io_dataOut_3777(dataOut[3777]),
.io_dataOut_3778(dataOut[3778]),
.io_dataOut_3779(dataOut[3779]),
.io_dataOut_3780(dataOut[3780]),
.io_dataOut_3781(dataOut[3781]),
.io_dataOut_3782(dataOut[3782]),
.io_dataOut_3783(dataOut[3783]),
.io_dataOut_3784(dataOut[3784]),
.io_dataOut_3785(dataOut[3785]),
.io_dataOut_3786(dataOut[3786]),
.io_dataOut_3787(dataOut[3787]),
.io_dataOut_3788(dataOut[3788]),
.io_dataOut_3789(dataOut[3789]),
.io_dataOut_3790(dataOut[3790]),
.io_dataOut_3791(dataOut[3791]),
.io_dataOut_3792(dataOut[3792]),
.io_dataOut_3793(dataOut[3793]),
.io_dataOut_3794(dataOut[3794]),
.io_dataOut_3795(dataOut[3795]),
.io_dataOut_3796(dataOut[3796]),
.io_dataOut_3797(dataOut[3797]),
.io_dataOut_3798(dataOut[3798]),
.io_dataOut_3799(dataOut[3799]),
.io_dataOut_3800(dataOut[3800]),
.io_dataOut_3801(dataOut[3801]),
.io_dataOut_3802(dataOut[3802]),
.io_dataOut_3803(dataOut[3803]),
.io_dataOut_3804(dataOut[3804]),
.io_dataOut_3805(dataOut[3805]),
.io_dataOut_3806(dataOut[3806]),
.io_dataOut_3807(dataOut[3807]),
.io_dataOut_3808(dataOut[3808]),
.io_dataOut_3809(dataOut[3809]),
.io_dataOut_3810(dataOut[3810]),
.io_dataOut_3811(dataOut[3811]),
.io_dataOut_3812(dataOut[3812]),
.io_dataOut_3813(dataOut[3813]),
.io_dataOut_3814(dataOut[3814]),
.io_dataOut_3815(dataOut[3815]),
.io_dataOut_3816(dataOut[3816]),
.io_dataOut_3817(dataOut[3817]),
.io_dataOut_3818(dataOut[3818]),
.io_dataOut_3819(dataOut[3819]),
.io_dataOut_3820(dataOut[3820]),
.io_dataOut_3821(dataOut[3821]),
.io_dataOut_3822(dataOut[3822]),
.io_dataOut_3823(dataOut[3823]),
.io_dataOut_3824(dataOut[3824]),
.io_dataOut_3825(dataOut[3825]),
.io_dataOut_3826(dataOut[3826]),
.io_dataOut_3827(dataOut[3827]),
.io_dataOut_3828(dataOut[3828]),
.io_dataOut_3829(dataOut[3829]),
.io_dataOut_3830(dataOut[3830]),
.io_dataOut_3831(dataOut[3831]),
.io_dataOut_3832(dataOut[3832]),
.io_dataOut_3833(dataOut[3833]),
.io_dataOut_3834(dataOut[3834]),
.io_dataOut_3835(dataOut[3835]),
.io_dataOut_3836(dataOut[3836]),
.io_dataOut_3837(dataOut[3837]),
.io_dataOut_3838(dataOut[3838]),
.io_dataOut_3839(dataOut[3839]),
.io_dataOut_3840(dataOut[3840]),
.io_dataOut_3841(dataOut[3841]),
.io_dataOut_3842(dataOut[3842]),
.io_dataOut_3843(dataOut[3843]),
.io_dataOut_3844(dataOut[3844]),
.io_dataOut_3845(dataOut[3845]),
.io_dataOut_3846(dataOut[3846]),
.io_dataOut_3847(dataOut[3847]),
.io_dataOut_3848(dataOut[3848]),
.io_dataOut_3849(dataOut[3849]),
.io_dataOut_3850(dataOut[3850]),
.io_dataOut_3851(dataOut[3851]),
.io_dataOut_3852(dataOut[3852]),
.io_dataOut_3853(dataOut[3853]),
.io_dataOut_3854(dataOut[3854]),
.io_dataOut_3855(dataOut[3855]),
.io_dataOut_3856(dataOut[3856]),
.io_dataOut_3857(dataOut[3857]),
.io_dataOut_3858(dataOut[3858]),
.io_dataOut_3859(dataOut[3859]),
.io_dataOut_3860(dataOut[3860]),
.io_dataOut_3861(dataOut[3861]),
.io_dataOut_3862(dataOut[3862]),
.io_dataOut_3863(dataOut[3863]),
.io_dataOut_3864(dataOut[3864]),
.io_dataOut_3865(dataOut[3865]),
.io_dataOut_3866(dataOut[3866]),
.io_dataOut_3867(dataOut[3867]),
.io_dataOut_3868(dataOut[3868]),
.io_dataOut_3869(dataOut[3869]),
.io_dataOut_3870(dataOut[3870]),
.io_dataOut_3871(dataOut[3871]),
.io_dataOut_3872(dataOut[3872]),
.io_dataOut_3873(dataOut[3873]),
.io_dataOut_3874(dataOut[3874]),
.io_dataOut_3875(dataOut[3875]),
.io_dataOut_3876(dataOut[3876]),
.io_dataOut_3877(dataOut[3877]),
.io_dataOut_3878(dataOut[3878]),
.io_dataOut_3879(dataOut[3879]),
.io_dataOut_3880(dataOut[3880]),
.io_dataOut_3881(dataOut[3881]),
.io_dataOut_3882(dataOut[3882]),
.io_dataOut_3883(dataOut[3883]),
.io_dataOut_3884(dataOut[3884]),
.io_dataOut_3885(dataOut[3885]),
.io_dataOut_3886(dataOut[3886]),
.io_dataOut_3887(dataOut[3887]),
.io_dataOut_3888(dataOut[3888]),
.io_dataOut_3889(dataOut[3889]),
.io_dataOut_3890(dataOut[3890]),
.io_dataOut_3891(dataOut[3891]),
.io_dataOut_3892(dataOut[3892]),
.io_dataOut_3893(dataOut[3893]),
.io_dataOut_3894(dataOut[3894]),
.io_dataOut_3895(dataOut[3895]),
.io_dataOut_3896(dataOut[3896]),
.io_dataOut_3897(dataOut[3897]),
.io_dataOut_3898(dataOut[3898]),
.io_dataOut_3899(dataOut[3899]),
.io_dataOut_3900(dataOut[3900]),
.io_dataOut_3901(dataOut[3901]),
.io_dataOut_3902(dataOut[3902]),
.io_dataOut_3903(dataOut[3903]),
.io_dataOut_3904(dataOut[3904]),
.io_dataOut_3905(dataOut[3905]),
.io_dataOut_3906(dataOut[3906]),
.io_dataOut_3907(dataOut[3907]),
.io_dataOut_3908(dataOut[3908]),
.io_dataOut_3909(dataOut[3909]),
.io_dataOut_3910(dataOut[3910]),
.io_dataOut_3911(dataOut[3911]),
.io_dataOut_3912(dataOut[3912]),
.io_dataOut_3913(dataOut[3913]),
.io_dataOut_3914(dataOut[3914]),
.io_dataOut_3915(dataOut[3915]),
.io_dataOut_3916(dataOut[3916]),
.io_dataOut_3917(dataOut[3917]),
.io_dataOut_3918(dataOut[3918]),
.io_dataOut_3919(dataOut[3919]),
.io_dataOut_3920(dataOut[3920]),
.io_dataOut_3921(dataOut[3921]),
.io_dataOut_3922(dataOut[3922]),
.io_dataOut_3923(dataOut[3923]),
.io_dataOut_3924(dataOut[3924]),
.io_dataOut_3925(dataOut[3925]),
.io_dataOut_3926(dataOut[3926]),
.io_dataOut_3927(dataOut[3927]),
.io_dataOut_3928(dataOut[3928]),
.io_dataOut_3929(dataOut[3929]),
.io_dataOut_3930(dataOut[3930]),
.io_dataOut_3931(dataOut[3931]),
.io_dataOut_3932(dataOut[3932]),
.io_dataOut_3933(dataOut[3933]),
.io_dataOut_3934(dataOut[3934]),
.io_dataOut_3935(dataOut[3935]),
.io_dataOut_3936(dataOut[3936]),
.io_dataOut_3937(dataOut[3937]),
.io_dataOut_3938(dataOut[3938]),
.io_dataOut_3939(dataOut[3939]),
.io_dataOut_3940(dataOut[3940]),
.io_dataOut_3941(dataOut[3941]),
.io_dataOut_3942(dataOut[3942]),
.io_dataOut_3943(dataOut[3943]),
.io_dataOut_3944(dataOut[3944]),
.io_dataOut_3945(dataOut[3945]),
.io_dataOut_3946(dataOut[3946]),
.io_dataOut_3947(dataOut[3947]),
.io_dataOut_3948(dataOut[3948]),
.io_dataOut_3949(dataOut[3949]),
.io_dataOut_3950(dataOut[3950]),
.io_dataOut_3951(dataOut[3951]),
.io_dataOut_3952(dataOut[3952]),
.io_dataOut_3953(dataOut[3953]),
.io_dataOut_3954(dataOut[3954]),
.io_dataOut_3955(dataOut[3955]),
.io_dataOut_3956(dataOut[3956]),
.io_dataOut_3957(dataOut[3957]),
.io_dataOut_3958(dataOut[3958]),
.io_dataOut_3959(dataOut[3959]),
.io_dataOut_3960(dataOut[3960]),
.io_dataOut_3961(dataOut[3961]),
.io_dataOut_3962(dataOut[3962]),
.io_dataOut_3963(dataOut[3963]),
.io_dataOut_3964(dataOut[3964]),
.io_dataOut_3965(dataOut[3965]),
.io_dataOut_3966(dataOut[3966]),
.io_dataOut_3967(dataOut[3967]),
.io_dataOut_3968(dataOut[3968]),
.io_dataOut_3969(dataOut[3969]),
.io_dataOut_3970(dataOut[3970]),
.io_dataOut_3971(dataOut[3971]),
.io_dataOut_3972(dataOut[3972]),
.io_dataOut_3973(dataOut[3973]),
.io_dataOut_3974(dataOut[3974]),
.io_dataOut_3975(dataOut[3975]),
.io_dataOut_3976(dataOut[3976]),
.io_dataOut_3977(dataOut[3977]),
.io_dataOut_3978(dataOut[3978]),
.io_dataOut_3979(dataOut[3979]),
.io_dataOut_3980(dataOut[3980]),
.io_dataOut_3981(dataOut[3981]),
.io_dataOut_3982(dataOut[3982]),
.io_dataOut_3983(dataOut[3983]),
.io_dataOut_3984(dataOut[3984]),
.io_dataOut_3985(dataOut[3985]),
.io_dataOut_3986(dataOut[3986]),
.io_dataOut_3987(dataOut[3987]),
.io_dataOut_3988(dataOut[3988]),
.io_dataOut_3989(dataOut[3989]),
.io_dataOut_3990(dataOut[3990]),
.io_dataOut_3991(dataOut[3991]),
.io_dataOut_3992(dataOut[3992]),
.io_dataOut_3993(dataOut[3993]),
.io_dataOut_3994(dataOut[3994]),
.io_dataOut_3995(dataOut[3995]),
.io_dataOut_3996(dataOut[3996]),
.io_dataOut_3997(dataOut[3997]),
.io_dataOut_3998(dataOut[3998]),
.io_dataOut_3999(dataOut[3999]),
.io_dataOut_4000(dataOut[4000]),
.io_dataOut_4001(dataOut[4001]),
.io_dataOut_4002(dataOut[4002]),
.io_dataOut_4003(dataOut[4003]),
.io_dataOut_4004(dataOut[4004]),
.io_dataOut_4005(dataOut[4005]),
.io_dataOut_4006(dataOut[4006]),
.io_dataOut_4007(dataOut[4007]),
.io_dataOut_4008(dataOut[4008]),
.io_dataOut_4009(dataOut[4009]),
.io_dataOut_4010(dataOut[4010]),
.io_dataOut_4011(dataOut[4011]),
.io_dataOut_4012(dataOut[4012]),
.io_dataOut_4013(dataOut[4013]),
.io_dataOut_4014(dataOut[4014]),
.io_dataOut_4015(dataOut[4015]),
.io_dataOut_4016(dataOut[4016]),
.io_dataOut_4017(dataOut[4017]),
.io_dataOut_4018(dataOut[4018]),
.io_dataOut_4019(dataOut[4019]),
.io_dataOut_4020(dataOut[4020]),
.io_dataOut_4021(dataOut[4021]),
.io_dataOut_4022(dataOut[4022]),
.io_dataOut_4023(dataOut[4023]),
.io_dataOut_4024(dataOut[4024]),
.io_dataOut_4025(dataOut[4025]),
.io_dataOut_4026(dataOut[4026]),
.io_dataOut_4027(dataOut[4027]),
.io_dataOut_4028(dataOut[4028]),
.io_dataOut_4029(dataOut[4029]),
.io_dataOut_4030(dataOut[4030]),
.io_dataOut_4031(dataOut[4031]),
.io_dataOut_4032(dataOut[4032]),
.io_dataOut_4033(dataOut[4033]),
.io_dataOut_4034(dataOut[4034]),
.io_dataOut_4035(dataOut[4035]),
.io_dataOut_4036(dataOut[4036]),
.io_dataOut_4037(dataOut[4037]),
.io_dataOut_4038(dataOut[4038]),
.io_dataOut_4039(dataOut[4039]),
.io_dataOut_4040(dataOut[4040]),
.io_dataOut_4041(dataOut[4041]),
.io_dataOut_4042(dataOut[4042]),
.io_dataOut_4043(dataOut[4043]),
.io_dataOut_4044(dataOut[4044]),
.io_dataOut_4045(dataOut[4045]),
.io_dataOut_4046(dataOut[4046]),
.io_dataOut_4047(dataOut[4047]),
.io_dataOut_4048(dataOut[4048]),
.io_dataOut_4049(dataOut[4049]),
.io_dataOut_4050(dataOut[4050]),
.io_dataOut_4051(dataOut[4051]),
.io_dataOut_4052(dataOut[4052]),
.io_dataOut_4053(dataOut[4053]),
.io_dataOut_4054(dataOut[4054]),
.io_dataOut_4055(dataOut[4055]),
.io_dataOut_4056(dataOut[4056]),
.io_dataOut_4057(dataOut[4057]),
.io_dataOut_4058(dataOut[4058]),
.io_dataOut_4059(dataOut[4059]),
.io_dataOut_4060(dataOut[4060]),
.io_dataOut_4061(dataOut[4061]),
.io_dataOut_4062(dataOut[4062]),
.io_dataOut_4063(dataOut[4063]),
.io_dataOut_4064(dataOut[4064]),
.io_dataOut_4065(dataOut[4065]),
.io_dataOut_4066(dataOut[4066]),
.io_dataOut_4067(dataOut[4067]),
.io_dataOut_4068(dataOut[4068]),
.io_dataOut_4069(dataOut[4069]),
.io_dataOut_4070(dataOut[4070]),
.io_dataOut_4071(dataOut[4071]),
.io_dataOut_4072(dataOut[4072]),
.io_dataOut_4073(dataOut[4073]),
.io_dataOut_4074(dataOut[4074]),
.io_dataOut_4075(dataOut[4075]),
.io_dataOut_4076(dataOut[4076]),
.io_dataOut_4077(dataOut[4077]),
.io_dataOut_4078(dataOut[4078]),
.io_dataOut_4079(dataOut[4079]),
.io_dataOut_4080(dataOut[4080]),
.io_dataOut_4081(dataOut[4081]),
.io_dataOut_4082(dataOut[4082]),
.io_dataOut_4083(dataOut[4083]),
.io_dataOut_4084(dataOut[4084]),
.io_dataOut_4085(dataOut[4085]),
.io_dataOut_4086(dataOut[4086]),
.io_dataOut_4087(dataOut[4087]),
.io_dataOut_4088(dataOut[4088]),
.io_dataOut_4089(dataOut[4089]),
.io_dataOut_4090(dataOut[4090]),
.io_dataOut_4091(dataOut[4091]),
.io_dataOut_4092(dataOut[4092]),
.io_dataOut_4093(dataOut[4093]),
.io_dataOut_4094(dataOut[4094]),
.io_dataOut_4095(dataOut[4095])
         );

endmodule

