// Wrapper for the toplevel module, which is the combination of the chisel
// implementation for the codeword generator and the compressorOutput

module lz77AndHuffmanWrapper(
         input clock,
         input reset,
         input [7:0] dataIn [0:4095],
         output [7:0] dataOut [0:4095],
         output matchingBytes [0:4095],
         output [12:0] numberOfMatchingBytes,
         output [12:0] lz77CompressedBytes,
         output [12:0] huffmanCompressedBytes,
         output finished
       );
       wire inValid, inReady, outReady, outValid;

lz77AndHuffman wrapped(
.clock(clock),
.reset(reset),
.io_finished(finished),
.io_in_0(dataIn[0]),
.io_in_1(dataIn[1]),
.io_in_2(dataIn[2]),
.io_in_3(dataIn[3]),
.io_in_4(dataIn[4]),
.io_in_5(dataIn[5]),
.io_in_6(dataIn[6]),
.io_in_7(dataIn[7]),
.io_in_8(dataIn[8]),
.io_in_9(dataIn[9]),
.io_in_10(dataIn[10]),
.io_in_11(dataIn[11]),
.io_in_12(dataIn[12]),
.io_in_13(dataIn[13]),
.io_in_14(dataIn[14]),
.io_in_15(dataIn[15]),
.io_in_16(dataIn[16]),
.io_in_17(dataIn[17]),
.io_in_18(dataIn[18]),
.io_in_19(dataIn[19]),
.io_in_20(dataIn[20]),
.io_in_21(dataIn[21]),
.io_in_22(dataIn[22]),
.io_in_23(dataIn[23]),
.io_in_24(dataIn[24]),
.io_in_25(dataIn[25]),
.io_in_26(dataIn[26]),
.io_in_27(dataIn[27]),
.io_in_28(dataIn[28]),
.io_in_29(dataIn[29]),
.io_in_30(dataIn[30]),
.io_in_31(dataIn[31]),
.io_in_32(dataIn[32]),
.io_in_33(dataIn[33]),
.io_in_34(dataIn[34]),
.io_in_35(dataIn[35]),
.io_in_36(dataIn[36]),
.io_in_37(dataIn[37]),
.io_in_38(dataIn[38]),
.io_in_39(dataIn[39]),
.io_in_40(dataIn[40]),
.io_in_41(dataIn[41]),
.io_in_42(dataIn[42]),
.io_in_43(dataIn[43]),
.io_in_44(dataIn[44]),
.io_in_45(dataIn[45]),
.io_in_46(dataIn[46]),
.io_in_47(dataIn[47]),
.io_in_48(dataIn[48]),
.io_in_49(dataIn[49]),
.io_in_50(dataIn[50]),
.io_in_51(dataIn[51]),
.io_in_52(dataIn[52]),
.io_in_53(dataIn[53]),
.io_in_54(dataIn[54]),
.io_in_55(dataIn[55]),
.io_in_56(dataIn[56]),
.io_in_57(dataIn[57]),
.io_in_58(dataIn[58]),
.io_in_59(dataIn[59]),
.io_in_60(dataIn[60]),
.io_in_61(dataIn[61]),
.io_in_62(dataIn[62]),
.io_in_63(dataIn[63]),
.io_in_64(dataIn[64]),
.io_in_65(dataIn[65]),
.io_in_66(dataIn[66]),
.io_in_67(dataIn[67]),
.io_in_68(dataIn[68]),
.io_in_69(dataIn[69]),
.io_in_70(dataIn[70]),
.io_in_71(dataIn[71]),
.io_in_72(dataIn[72]),
.io_in_73(dataIn[73]),
.io_in_74(dataIn[74]),
.io_in_75(dataIn[75]),
.io_in_76(dataIn[76]),
.io_in_77(dataIn[77]),
.io_in_78(dataIn[78]),
.io_in_79(dataIn[79]),
.io_in_80(dataIn[80]),
.io_in_81(dataIn[81]),
.io_in_82(dataIn[82]),
.io_in_83(dataIn[83]),
.io_in_84(dataIn[84]),
.io_in_85(dataIn[85]),
.io_in_86(dataIn[86]),
.io_in_87(dataIn[87]),
.io_in_88(dataIn[88]),
.io_in_89(dataIn[89]),
.io_in_90(dataIn[90]),
.io_in_91(dataIn[91]),
.io_in_92(dataIn[92]),
.io_in_93(dataIn[93]),
.io_in_94(dataIn[94]),
.io_in_95(dataIn[95]),
.io_in_96(dataIn[96]),
.io_in_97(dataIn[97]),
.io_in_98(dataIn[98]),
.io_in_99(dataIn[99]),
.io_in_100(dataIn[100]),
.io_in_101(dataIn[101]),
.io_in_102(dataIn[102]),
.io_in_103(dataIn[103]),
.io_in_104(dataIn[104]),
.io_in_105(dataIn[105]),
.io_in_106(dataIn[106]),
.io_in_107(dataIn[107]),
.io_in_108(dataIn[108]),
.io_in_109(dataIn[109]),
.io_in_110(dataIn[110]),
.io_in_111(dataIn[111]),
.io_in_112(dataIn[112]),
.io_in_113(dataIn[113]),
.io_in_114(dataIn[114]),
.io_in_115(dataIn[115]),
.io_in_116(dataIn[116]),
.io_in_117(dataIn[117]),
.io_in_118(dataIn[118]),
.io_in_119(dataIn[119]),
.io_in_120(dataIn[120]),
.io_in_121(dataIn[121]),
.io_in_122(dataIn[122]),
.io_in_123(dataIn[123]),
.io_in_124(dataIn[124]),
.io_in_125(dataIn[125]),
.io_in_126(dataIn[126]),
.io_in_127(dataIn[127]),
.io_in_128(dataIn[128]),
.io_in_129(dataIn[129]),
.io_in_130(dataIn[130]),
.io_in_131(dataIn[131]),
.io_in_132(dataIn[132]),
.io_in_133(dataIn[133]),
.io_in_134(dataIn[134]),
.io_in_135(dataIn[135]),
.io_in_136(dataIn[136]),
.io_in_137(dataIn[137]),
.io_in_138(dataIn[138]),
.io_in_139(dataIn[139]),
.io_in_140(dataIn[140]),
.io_in_141(dataIn[141]),
.io_in_142(dataIn[142]),
.io_in_143(dataIn[143]),
.io_in_144(dataIn[144]),
.io_in_145(dataIn[145]),
.io_in_146(dataIn[146]),
.io_in_147(dataIn[147]),
.io_in_148(dataIn[148]),
.io_in_149(dataIn[149]),
.io_in_150(dataIn[150]),
.io_in_151(dataIn[151]),
.io_in_152(dataIn[152]),
.io_in_153(dataIn[153]),
.io_in_154(dataIn[154]),
.io_in_155(dataIn[155]),
.io_in_156(dataIn[156]),
.io_in_157(dataIn[157]),
.io_in_158(dataIn[158]),
.io_in_159(dataIn[159]),
.io_in_160(dataIn[160]),
.io_in_161(dataIn[161]),
.io_in_162(dataIn[162]),
.io_in_163(dataIn[163]),
.io_in_164(dataIn[164]),
.io_in_165(dataIn[165]),
.io_in_166(dataIn[166]),
.io_in_167(dataIn[167]),
.io_in_168(dataIn[168]),
.io_in_169(dataIn[169]),
.io_in_170(dataIn[170]),
.io_in_171(dataIn[171]),
.io_in_172(dataIn[172]),
.io_in_173(dataIn[173]),
.io_in_174(dataIn[174]),
.io_in_175(dataIn[175]),
.io_in_176(dataIn[176]),
.io_in_177(dataIn[177]),
.io_in_178(dataIn[178]),
.io_in_179(dataIn[179]),
.io_in_180(dataIn[180]),
.io_in_181(dataIn[181]),
.io_in_182(dataIn[182]),
.io_in_183(dataIn[183]),
.io_in_184(dataIn[184]),
.io_in_185(dataIn[185]),
.io_in_186(dataIn[186]),
.io_in_187(dataIn[187]),
.io_in_188(dataIn[188]),
.io_in_189(dataIn[189]),
.io_in_190(dataIn[190]),
.io_in_191(dataIn[191]),
.io_in_192(dataIn[192]),
.io_in_193(dataIn[193]),
.io_in_194(dataIn[194]),
.io_in_195(dataIn[195]),
.io_in_196(dataIn[196]),
.io_in_197(dataIn[197]),
.io_in_198(dataIn[198]),
.io_in_199(dataIn[199]),
.io_in_200(dataIn[200]),
.io_in_201(dataIn[201]),
.io_in_202(dataIn[202]),
.io_in_203(dataIn[203]),
.io_in_204(dataIn[204]),
.io_in_205(dataIn[205]),
.io_in_206(dataIn[206]),
.io_in_207(dataIn[207]),
.io_in_208(dataIn[208]),
.io_in_209(dataIn[209]),
.io_in_210(dataIn[210]),
.io_in_211(dataIn[211]),
.io_in_212(dataIn[212]),
.io_in_213(dataIn[213]),
.io_in_214(dataIn[214]),
.io_in_215(dataIn[215]),
.io_in_216(dataIn[216]),
.io_in_217(dataIn[217]),
.io_in_218(dataIn[218]),
.io_in_219(dataIn[219]),
.io_in_220(dataIn[220]),
.io_in_221(dataIn[221]),
.io_in_222(dataIn[222]),
.io_in_223(dataIn[223]),
.io_in_224(dataIn[224]),
.io_in_225(dataIn[225]),
.io_in_226(dataIn[226]),
.io_in_227(dataIn[227]),
.io_in_228(dataIn[228]),
.io_in_229(dataIn[229]),
.io_in_230(dataIn[230]),
.io_in_231(dataIn[231]),
.io_in_232(dataIn[232]),
.io_in_233(dataIn[233]),
.io_in_234(dataIn[234]),
.io_in_235(dataIn[235]),
.io_in_236(dataIn[236]),
.io_in_237(dataIn[237]),
.io_in_238(dataIn[238]),
.io_in_239(dataIn[239]),
.io_in_240(dataIn[240]),
.io_in_241(dataIn[241]),
.io_in_242(dataIn[242]),
.io_in_243(dataIn[243]),
.io_in_244(dataIn[244]),
.io_in_245(dataIn[245]),
.io_in_246(dataIn[246]),
.io_in_247(dataIn[247]),
.io_in_248(dataIn[248]),
.io_in_249(dataIn[249]),
.io_in_250(dataIn[250]),
.io_in_251(dataIn[251]),
.io_in_252(dataIn[252]),
.io_in_253(dataIn[253]),
.io_in_254(dataIn[254]),
.io_in_255(dataIn[255]),
.io_in_256(dataIn[256]),
.io_in_257(dataIn[257]),
.io_in_258(dataIn[258]),
.io_in_259(dataIn[259]),
.io_in_260(dataIn[260]),
.io_in_261(dataIn[261]),
.io_in_262(dataIn[262]),
.io_in_263(dataIn[263]),
.io_in_264(dataIn[264]),
.io_in_265(dataIn[265]),
.io_in_266(dataIn[266]),
.io_in_267(dataIn[267]),
.io_in_268(dataIn[268]),
.io_in_269(dataIn[269]),
.io_in_270(dataIn[270]),
.io_in_271(dataIn[271]),
.io_in_272(dataIn[272]),
.io_in_273(dataIn[273]),
.io_in_274(dataIn[274]),
.io_in_275(dataIn[275]),
.io_in_276(dataIn[276]),
.io_in_277(dataIn[277]),
.io_in_278(dataIn[278]),
.io_in_279(dataIn[279]),
.io_in_280(dataIn[280]),
.io_in_281(dataIn[281]),
.io_in_282(dataIn[282]),
.io_in_283(dataIn[283]),
.io_in_284(dataIn[284]),
.io_in_285(dataIn[285]),
.io_in_286(dataIn[286]),
.io_in_287(dataIn[287]),
.io_in_288(dataIn[288]),
.io_in_289(dataIn[289]),
.io_in_290(dataIn[290]),
.io_in_291(dataIn[291]),
.io_in_292(dataIn[292]),
.io_in_293(dataIn[293]),
.io_in_294(dataIn[294]),
.io_in_295(dataIn[295]),
.io_in_296(dataIn[296]),
.io_in_297(dataIn[297]),
.io_in_298(dataIn[298]),
.io_in_299(dataIn[299]),
.io_in_300(dataIn[300]),
.io_in_301(dataIn[301]),
.io_in_302(dataIn[302]),
.io_in_303(dataIn[303]),
.io_in_304(dataIn[304]),
.io_in_305(dataIn[305]),
.io_in_306(dataIn[306]),
.io_in_307(dataIn[307]),
.io_in_308(dataIn[308]),
.io_in_309(dataIn[309]),
.io_in_310(dataIn[310]),
.io_in_311(dataIn[311]),
.io_in_312(dataIn[312]),
.io_in_313(dataIn[313]),
.io_in_314(dataIn[314]),
.io_in_315(dataIn[315]),
.io_in_316(dataIn[316]),
.io_in_317(dataIn[317]),
.io_in_318(dataIn[318]),
.io_in_319(dataIn[319]),
.io_in_320(dataIn[320]),
.io_in_321(dataIn[321]),
.io_in_322(dataIn[322]),
.io_in_323(dataIn[323]),
.io_in_324(dataIn[324]),
.io_in_325(dataIn[325]),
.io_in_326(dataIn[326]),
.io_in_327(dataIn[327]),
.io_in_328(dataIn[328]),
.io_in_329(dataIn[329]),
.io_in_330(dataIn[330]),
.io_in_331(dataIn[331]),
.io_in_332(dataIn[332]),
.io_in_333(dataIn[333]),
.io_in_334(dataIn[334]),
.io_in_335(dataIn[335]),
.io_in_336(dataIn[336]),
.io_in_337(dataIn[337]),
.io_in_338(dataIn[338]),
.io_in_339(dataIn[339]),
.io_in_340(dataIn[340]),
.io_in_341(dataIn[341]),
.io_in_342(dataIn[342]),
.io_in_343(dataIn[343]),
.io_in_344(dataIn[344]),
.io_in_345(dataIn[345]),
.io_in_346(dataIn[346]),
.io_in_347(dataIn[347]),
.io_in_348(dataIn[348]),
.io_in_349(dataIn[349]),
.io_in_350(dataIn[350]),
.io_in_351(dataIn[351]),
.io_in_352(dataIn[352]),
.io_in_353(dataIn[353]),
.io_in_354(dataIn[354]),
.io_in_355(dataIn[355]),
.io_in_356(dataIn[356]),
.io_in_357(dataIn[357]),
.io_in_358(dataIn[358]),
.io_in_359(dataIn[359]),
.io_in_360(dataIn[360]),
.io_in_361(dataIn[361]),
.io_in_362(dataIn[362]),
.io_in_363(dataIn[363]),
.io_in_364(dataIn[364]),
.io_in_365(dataIn[365]),
.io_in_366(dataIn[366]),
.io_in_367(dataIn[367]),
.io_in_368(dataIn[368]),
.io_in_369(dataIn[369]),
.io_in_370(dataIn[370]),
.io_in_371(dataIn[371]),
.io_in_372(dataIn[372]),
.io_in_373(dataIn[373]),
.io_in_374(dataIn[374]),
.io_in_375(dataIn[375]),
.io_in_376(dataIn[376]),
.io_in_377(dataIn[377]),
.io_in_378(dataIn[378]),
.io_in_379(dataIn[379]),
.io_in_380(dataIn[380]),
.io_in_381(dataIn[381]),
.io_in_382(dataIn[382]),
.io_in_383(dataIn[383]),
.io_in_384(dataIn[384]),
.io_in_385(dataIn[385]),
.io_in_386(dataIn[386]),
.io_in_387(dataIn[387]),
.io_in_388(dataIn[388]),
.io_in_389(dataIn[389]),
.io_in_390(dataIn[390]),
.io_in_391(dataIn[391]),
.io_in_392(dataIn[392]),
.io_in_393(dataIn[393]),
.io_in_394(dataIn[394]),
.io_in_395(dataIn[395]),
.io_in_396(dataIn[396]),
.io_in_397(dataIn[397]),
.io_in_398(dataIn[398]),
.io_in_399(dataIn[399]),
.io_in_400(dataIn[400]),
.io_in_401(dataIn[401]),
.io_in_402(dataIn[402]),
.io_in_403(dataIn[403]),
.io_in_404(dataIn[404]),
.io_in_405(dataIn[405]),
.io_in_406(dataIn[406]),
.io_in_407(dataIn[407]),
.io_in_408(dataIn[408]),
.io_in_409(dataIn[409]),
.io_in_410(dataIn[410]),
.io_in_411(dataIn[411]),
.io_in_412(dataIn[412]),
.io_in_413(dataIn[413]),
.io_in_414(dataIn[414]),
.io_in_415(dataIn[415]),
.io_in_416(dataIn[416]),
.io_in_417(dataIn[417]),
.io_in_418(dataIn[418]),
.io_in_419(dataIn[419]),
.io_in_420(dataIn[420]),
.io_in_421(dataIn[421]),
.io_in_422(dataIn[422]),
.io_in_423(dataIn[423]),
.io_in_424(dataIn[424]),
.io_in_425(dataIn[425]),
.io_in_426(dataIn[426]),
.io_in_427(dataIn[427]),
.io_in_428(dataIn[428]),
.io_in_429(dataIn[429]),
.io_in_430(dataIn[430]),
.io_in_431(dataIn[431]),
.io_in_432(dataIn[432]),
.io_in_433(dataIn[433]),
.io_in_434(dataIn[434]),
.io_in_435(dataIn[435]),
.io_in_436(dataIn[436]),
.io_in_437(dataIn[437]),
.io_in_438(dataIn[438]),
.io_in_439(dataIn[439]),
.io_in_440(dataIn[440]),
.io_in_441(dataIn[441]),
.io_in_442(dataIn[442]),
.io_in_443(dataIn[443]),
.io_in_444(dataIn[444]),
.io_in_445(dataIn[445]),
.io_in_446(dataIn[446]),
.io_in_447(dataIn[447]),
.io_in_448(dataIn[448]),
.io_in_449(dataIn[449]),
.io_in_450(dataIn[450]),
.io_in_451(dataIn[451]),
.io_in_452(dataIn[452]),
.io_in_453(dataIn[453]),
.io_in_454(dataIn[454]),
.io_in_455(dataIn[455]),
.io_in_456(dataIn[456]),
.io_in_457(dataIn[457]),
.io_in_458(dataIn[458]),
.io_in_459(dataIn[459]),
.io_in_460(dataIn[460]),
.io_in_461(dataIn[461]),
.io_in_462(dataIn[462]),
.io_in_463(dataIn[463]),
.io_in_464(dataIn[464]),
.io_in_465(dataIn[465]),
.io_in_466(dataIn[466]),
.io_in_467(dataIn[467]),
.io_in_468(dataIn[468]),
.io_in_469(dataIn[469]),
.io_in_470(dataIn[470]),
.io_in_471(dataIn[471]),
.io_in_472(dataIn[472]),
.io_in_473(dataIn[473]),
.io_in_474(dataIn[474]),
.io_in_475(dataIn[475]),
.io_in_476(dataIn[476]),
.io_in_477(dataIn[477]),
.io_in_478(dataIn[478]),
.io_in_479(dataIn[479]),
.io_in_480(dataIn[480]),
.io_in_481(dataIn[481]),
.io_in_482(dataIn[482]),
.io_in_483(dataIn[483]),
.io_in_484(dataIn[484]),
.io_in_485(dataIn[485]),
.io_in_486(dataIn[486]),
.io_in_487(dataIn[487]),
.io_in_488(dataIn[488]),
.io_in_489(dataIn[489]),
.io_in_490(dataIn[490]),
.io_in_491(dataIn[491]),
.io_in_492(dataIn[492]),
.io_in_493(dataIn[493]),
.io_in_494(dataIn[494]),
.io_in_495(dataIn[495]),
.io_in_496(dataIn[496]),
.io_in_497(dataIn[497]),
.io_in_498(dataIn[498]),
.io_in_499(dataIn[499]),
.io_in_500(dataIn[500]),
.io_in_501(dataIn[501]),
.io_in_502(dataIn[502]),
.io_in_503(dataIn[503]),
.io_in_504(dataIn[504]),
.io_in_505(dataIn[505]),
.io_in_506(dataIn[506]),
.io_in_507(dataIn[507]),
.io_in_508(dataIn[508]),
.io_in_509(dataIn[509]),
.io_in_510(dataIn[510]),
.io_in_511(dataIn[511]),
.io_in_512(dataIn[512]),
.io_in_513(dataIn[513]),
.io_in_514(dataIn[514]),
.io_in_515(dataIn[515]),
.io_in_516(dataIn[516]),
.io_in_517(dataIn[517]),
.io_in_518(dataIn[518]),
.io_in_519(dataIn[519]),
.io_in_520(dataIn[520]),
.io_in_521(dataIn[521]),
.io_in_522(dataIn[522]),
.io_in_523(dataIn[523]),
.io_in_524(dataIn[524]),
.io_in_525(dataIn[525]),
.io_in_526(dataIn[526]),
.io_in_527(dataIn[527]),
.io_in_528(dataIn[528]),
.io_in_529(dataIn[529]),
.io_in_530(dataIn[530]),
.io_in_531(dataIn[531]),
.io_in_532(dataIn[532]),
.io_in_533(dataIn[533]),
.io_in_534(dataIn[534]),
.io_in_535(dataIn[535]),
.io_in_536(dataIn[536]),
.io_in_537(dataIn[537]),
.io_in_538(dataIn[538]),
.io_in_539(dataIn[539]),
.io_in_540(dataIn[540]),
.io_in_541(dataIn[541]),
.io_in_542(dataIn[542]),
.io_in_543(dataIn[543]),
.io_in_544(dataIn[544]),
.io_in_545(dataIn[545]),
.io_in_546(dataIn[546]),
.io_in_547(dataIn[547]),
.io_in_548(dataIn[548]),
.io_in_549(dataIn[549]),
.io_in_550(dataIn[550]),
.io_in_551(dataIn[551]),
.io_in_552(dataIn[552]),
.io_in_553(dataIn[553]),
.io_in_554(dataIn[554]),
.io_in_555(dataIn[555]),
.io_in_556(dataIn[556]),
.io_in_557(dataIn[557]),
.io_in_558(dataIn[558]),
.io_in_559(dataIn[559]),
.io_in_560(dataIn[560]),
.io_in_561(dataIn[561]),
.io_in_562(dataIn[562]),
.io_in_563(dataIn[563]),
.io_in_564(dataIn[564]),
.io_in_565(dataIn[565]),
.io_in_566(dataIn[566]),
.io_in_567(dataIn[567]),
.io_in_568(dataIn[568]),
.io_in_569(dataIn[569]),
.io_in_570(dataIn[570]),
.io_in_571(dataIn[571]),
.io_in_572(dataIn[572]),
.io_in_573(dataIn[573]),
.io_in_574(dataIn[574]),
.io_in_575(dataIn[575]),
.io_in_576(dataIn[576]),
.io_in_577(dataIn[577]),
.io_in_578(dataIn[578]),
.io_in_579(dataIn[579]),
.io_in_580(dataIn[580]),
.io_in_581(dataIn[581]),
.io_in_582(dataIn[582]),
.io_in_583(dataIn[583]),
.io_in_584(dataIn[584]),
.io_in_585(dataIn[585]),
.io_in_586(dataIn[586]),
.io_in_587(dataIn[587]),
.io_in_588(dataIn[588]),
.io_in_589(dataIn[589]),
.io_in_590(dataIn[590]),
.io_in_591(dataIn[591]),
.io_in_592(dataIn[592]),
.io_in_593(dataIn[593]),
.io_in_594(dataIn[594]),
.io_in_595(dataIn[595]),
.io_in_596(dataIn[596]),
.io_in_597(dataIn[597]),
.io_in_598(dataIn[598]),
.io_in_599(dataIn[599]),
.io_in_600(dataIn[600]),
.io_in_601(dataIn[601]),
.io_in_602(dataIn[602]),
.io_in_603(dataIn[603]),
.io_in_604(dataIn[604]),
.io_in_605(dataIn[605]),
.io_in_606(dataIn[606]),
.io_in_607(dataIn[607]),
.io_in_608(dataIn[608]),
.io_in_609(dataIn[609]),
.io_in_610(dataIn[610]),
.io_in_611(dataIn[611]),
.io_in_612(dataIn[612]),
.io_in_613(dataIn[613]),
.io_in_614(dataIn[614]),
.io_in_615(dataIn[615]),
.io_in_616(dataIn[616]),
.io_in_617(dataIn[617]),
.io_in_618(dataIn[618]),
.io_in_619(dataIn[619]),
.io_in_620(dataIn[620]),
.io_in_621(dataIn[621]),
.io_in_622(dataIn[622]),
.io_in_623(dataIn[623]),
.io_in_624(dataIn[624]),
.io_in_625(dataIn[625]),
.io_in_626(dataIn[626]),
.io_in_627(dataIn[627]),
.io_in_628(dataIn[628]),
.io_in_629(dataIn[629]),
.io_in_630(dataIn[630]),
.io_in_631(dataIn[631]),
.io_in_632(dataIn[632]),
.io_in_633(dataIn[633]),
.io_in_634(dataIn[634]),
.io_in_635(dataIn[635]),
.io_in_636(dataIn[636]),
.io_in_637(dataIn[637]),
.io_in_638(dataIn[638]),
.io_in_639(dataIn[639]),
.io_in_640(dataIn[640]),
.io_in_641(dataIn[641]),
.io_in_642(dataIn[642]),
.io_in_643(dataIn[643]),
.io_in_644(dataIn[644]),
.io_in_645(dataIn[645]),
.io_in_646(dataIn[646]),
.io_in_647(dataIn[647]),
.io_in_648(dataIn[648]),
.io_in_649(dataIn[649]),
.io_in_650(dataIn[650]),
.io_in_651(dataIn[651]),
.io_in_652(dataIn[652]),
.io_in_653(dataIn[653]),
.io_in_654(dataIn[654]),
.io_in_655(dataIn[655]),
.io_in_656(dataIn[656]),
.io_in_657(dataIn[657]),
.io_in_658(dataIn[658]),
.io_in_659(dataIn[659]),
.io_in_660(dataIn[660]),
.io_in_661(dataIn[661]),
.io_in_662(dataIn[662]),
.io_in_663(dataIn[663]),
.io_in_664(dataIn[664]),
.io_in_665(dataIn[665]),
.io_in_666(dataIn[666]),
.io_in_667(dataIn[667]),
.io_in_668(dataIn[668]),
.io_in_669(dataIn[669]),
.io_in_670(dataIn[670]),
.io_in_671(dataIn[671]),
.io_in_672(dataIn[672]),
.io_in_673(dataIn[673]),
.io_in_674(dataIn[674]),
.io_in_675(dataIn[675]),
.io_in_676(dataIn[676]),
.io_in_677(dataIn[677]),
.io_in_678(dataIn[678]),
.io_in_679(dataIn[679]),
.io_in_680(dataIn[680]),
.io_in_681(dataIn[681]),
.io_in_682(dataIn[682]),
.io_in_683(dataIn[683]),
.io_in_684(dataIn[684]),
.io_in_685(dataIn[685]),
.io_in_686(dataIn[686]),
.io_in_687(dataIn[687]),
.io_in_688(dataIn[688]),
.io_in_689(dataIn[689]),
.io_in_690(dataIn[690]),
.io_in_691(dataIn[691]),
.io_in_692(dataIn[692]),
.io_in_693(dataIn[693]),
.io_in_694(dataIn[694]),
.io_in_695(dataIn[695]),
.io_in_696(dataIn[696]),
.io_in_697(dataIn[697]),
.io_in_698(dataIn[698]),
.io_in_699(dataIn[699]),
.io_in_700(dataIn[700]),
.io_in_701(dataIn[701]),
.io_in_702(dataIn[702]),
.io_in_703(dataIn[703]),
.io_in_704(dataIn[704]),
.io_in_705(dataIn[705]),
.io_in_706(dataIn[706]),
.io_in_707(dataIn[707]),
.io_in_708(dataIn[708]),
.io_in_709(dataIn[709]),
.io_in_710(dataIn[710]),
.io_in_711(dataIn[711]),
.io_in_712(dataIn[712]),
.io_in_713(dataIn[713]),
.io_in_714(dataIn[714]),
.io_in_715(dataIn[715]),
.io_in_716(dataIn[716]),
.io_in_717(dataIn[717]),
.io_in_718(dataIn[718]),
.io_in_719(dataIn[719]),
.io_in_720(dataIn[720]),
.io_in_721(dataIn[721]),
.io_in_722(dataIn[722]),
.io_in_723(dataIn[723]),
.io_in_724(dataIn[724]),
.io_in_725(dataIn[725]),
.io_in_726(dataIn[726]),
.io_in_727(dataIn[727]),
.io_in_728(dataIn[728]),
.io_in_729(dataIn[729]),
.io_in_730(dataIn[730]),
.io_in_731(dataIn[731]),
.io_in_732(dataIn[732]),
.io_in_733(dataIn[733]),
.io_in_734(dataIn[734]),
.io_in_735(dataIn[735]),
.io_in_736(dataIn[736]),
.io_in_737(dataIn[737]),
.io_in_738(dataIn[738]),
.io_in_739(dataIn[739]),
.io_in_740(dataIn[740]),
.io_in_741(dataIn[741]),
.io_in_742(dataIn[742]),
.io_in_743(dataIn[743]),
.io_in_744(dataIn[744]),
.io_in_745(dataIn[745]),
.io_in_746(dataIn[746]),
.io_in_747(dataIn[747]),
.io_in_748(dataIn[748]),
.io_in_749(dataIn[749]),
.io_in_750(dataIn[750]),
.io_in_751(dataIn[751]),
.io_in_752(dataIn[752]),
.io_in_753(dataIn[753]),
.io_in_754(dataIn[754]),
.io_in_755(dataIn[755]),
.io_in_756(dataIn[756]),
.io_in_757(dataIn[757]),
.io_in_758(dataIn[758]),
.io_in_759(dataIn[759]),
.io_in_760(dataIn[760]),
.io_in_761(dataIn[761]),
.io_in_762(dataIn[762]),
.io_in_763(dataIn[763]),
.io_in_764(dataIn[764]),
.io_in_765(dataIn[765]),
.io_in_766(dataIn[766]),
.io_in_767(dataIn[767]),
.io_in_768(dataIn[768]),
.io_in_769(dataIn[769]),
.io_in_770(dataIn[770]),
.io_in_771(dataIn[771]),
.io_in_772(dataIn[772]),
.io_in_773(dataIn[773]),
.io_in_774(dataIn[774]),
.io_in_775(dataIn[775]),
.io_in_776(dataIn[776]),
.io_in_777(dataIn[777]),
.io_in_778(dataIn[778]),
.io_in_779(dataIn[779]),
.io_in_780(dataIn[780]),
.io_in_781(dataIn[781]),
.io_in_782(dataIn[782]),
.io_in_783(dataIn[783]),
.io_in_784(dataIn[784]),
.io_in_785(dataIn[785]),
.io_in_786(dataIn[786]),
.io_in_787(dataIn[787]),
.io_in_788(dataIn[788]),
.io_in_789(dataIn[789]),
.io_in_790(dataIn[790]),
.io_in_791(dataIn[791]),
.io_in_792(dataIn[792]),
.io_in_793(dataIn[793]),
.io_in_794(dataIn[794]),
.io_in_795(dataIn[795]),
.io_in_796(dataIn[796]),
.io_in_797(dataIn[797]),
.io_in_798(dataIn[798]),
.io_in_799(dataIn[799]),
.io_in_800(dataIn[800]),
.io_in_801(dataIn[801]),
.io_in_802(dataIn[802]),
.io_in_803(dataIn[803]),
.io_in_804(dataIn[804]),
.io_in_805(dataIn[805]),
.io_in_806(dataIn[806]),
.io_in_807(dataIn[807]),
.io_in_808(dataIn[808]),
.io_in_809(dataIn[809]),
.io_in_810(dataIn[810]),
.io_in_811(dataIn[811]),
.io_in_812(dataIn[812]),
.io_in_813(dataIn[813]),
.io_in_814(dataIn[814]),
.io_in_815(dataIn[815]),
.io_in_816(dataIn[816]),
.io_in_817(dataIn[817]),
.io_in_818(dataIn[818]),
.io_in_819(dataIn[819]),
.io_in_820(dataIn[820]),
.io_in_821(dataIn[821]),
.io_in_822(dataIn[822]),
.io_in_823(dataIn[823]),
.io_in_824(dataIn[824]),
.io_in_825(dataIn[825]),
.io_in_826(dataIn[826]),
.io_in_827(dataIn[827]),
.io_in_828(dataIn[828]),
.io_in_829(dataIn[829]),
.io_in_830(dataIn[830]),
.io_in_831(dataIn[831]),
.io_in_832(dataIn[832]),
.io_in_833(dataIn[833]),
.io_in_834(dataIn[834]),
.io_in_835(dataIn[835]),
.io_in_836(dataIn[836]),
.io_in_837(dataIn[837]),
.io_in_838(dataIn[838]),
.io_in_839(dataIn[839]),
.io_in_840(dataIn[840]),
.io_in_841(dataIn[841]),
.io_in_842(dataIn[842]),
.io_in_843(dataIn[843]),
.io_in_844(dataIn[844]),
.io_in_845(dataIn[845]),
.io_in_846(dataIn[846]),
.io_in_847(dataIn[847]),
.io_in_848(dataIn[848]),
.io_in_849(dataIn[849]),
.io_in_850(dataIn[850]),
.io_in_851(dataIn[851]),
.io_in_852(dataIn[852]),
.io_in_853(dataIn[853]),
.io_in_854(dataIn[854]),
.io_in_855(dataIn[855]),
.io_in_856(dataIn[856]),
.io_in_857(dataIn[857]),
.io_in_858(dataIn[858]),
.io_in_859(dataIn[859]),
.io_in_860(dataIn[860]),
.io_in_861(dataIn[861]),
.io_in_862(dataIn[862]),
.io_in_863(dataIn[863]),
.io_in_864(dataIn[864]),
.io_in_865(dataIn[865]),
.io_in_866(dataIn[866]),
.io_in_867(dataIn[867]),
.io_in_868(dataIn[868]),
.io_in_869(dataIn[869]),
.io_in_870(dataIn[870]),
.io_in_871(dataIn[871]),
.io_in_872(dataIn[872]),
.io_in_873(dataIn[873]),
.io_in_874(dataIn[874]),
.io_in_875(dataIn[875]),
.io_in_876(dataIn[876]),
.io_in_877(dataIn[877]),
.io_in_878(dataIn[878]),
.io_in_879(dataIn[879]),
.io_in_880(dataIn[880]),
.io_in_881(dataIn[881]),
.io_in_882(dataIn[882]),
.io_in_883(dataIn[883]),
.io_in_884(dataIn[884]),
.io_in_885(dataIn[885]),
.io_in_886(dataIn[886]),
.io_in_887(dataIn[887]),
.io_in_888(dataIn[888]),
.io_in_889(dataIn[889]),
.io_in_890(dataIn[890]),
.io_in_891(dataIn[891]),
.io_in_892(dataIn[892]),
.io_in_893(dataIn[893]),
.io_in_894(dataIn[894]),
.io_in_895(dataIn[895]),
.io_in_896(dataIn[896]),
.io_in_897(dataIn[897]),
.io_in_898(dataIn[898]),
.io_in_899(dataIn[899]),
.io_in_900(dataIn[900]),
.io_in_901(dataIn[901]),
.io_in_902(dataIn[902]),
.io_in_903(dataIn[903]),
.io_in_904(dataIn[904]),
.io_in_905(dataIn[905]),
.io_in_906(dataIn[906]),
.io_in_907(dataIn[907]),
.io_in_908(dataIn[908]),
.io_in_909(dataIn[909]),
.io_in_910(dataIn[910]),
.io_in_911(dataIn[911]),
.io_in_912(dataIn[912]),
.io_in_913(dataIn[913]),
.io_in_914(dataIn[914]),
.io_in_915(dataIn[915]),
.io_in_916(dataIn[916]),
.io_in_917(dataIn[917]),
.io_in_918(dataIn[918]),
.io_in_919(dataIn[919]),
.io_in_920(dataIn[920]),
.io_in_921(dataIn[921]),
.io_in_922(dataIn[922]),
.io_in_923(dataIn[923]),
.io_in_924(dataIn[924]),
.io_in_925(dataIn[925]),
.io_in_926(dataIn[926]),
.io_in_927(dataIn[927]),
.io_in_928(dataIn[928]),
.io_in_929(dataIn[929]),
.io_in_930(dataIn[930]),
.io_in_931(dataIn[931]),
.io_in_932(dataIn[932]),
.io_in_933(dataIn[933]),
.io_in_934(dataIn[934]),
.io_in_935(dataIn[935]),
.io_in_936(dataIn[936]),
.io_in_937(dataIn[937]),
.io_in_938(dataIn[938]),
.io_in_939(dataIn[939]),
.io_in_940(dataIn[940]),
.io_in_941(dataIn[941]),
.io_in_942(dataIn[942]),
.io_in_943(dataIn[943]),
.io_in_944(dataIn[944]),
.io_in_945(dataIn[945]),
.io_in_946(dataIn[946]),
.io_in_947(dataIn[947]),
.io_in_948(dataIn[948]),
.io_in_949(dataIn[949]),
.io_in_950(dataIn[950]),
.io_in_951(dataIn[951]),
.io_in_952(dataIn[952]),
.io_in_953(dataIn[953]),
.io_in_954(dataIn[954]),
.io_in_955(dataIn[955]),
.io_in_956(dataIn[956]),
.io_in_957(dataIn[957]),
.io_in_958(dataIn[958]),
.io_in_959(dataIn[959]),
.io_in_960(dataIn[960]),
.io_in_961(dataIn[961]),
.io_in_962(dataIn[962]),
.io_in_963(dataIn[963]),
.io_in_964(dataIn[964]),
.io_in_965(dataIn[965]),
.io_in_966(dataIn[966]),
.io_in_967(dataIn[967]),
.io_in_968(dataIn[968]),
.io_in_969(dataIn[969]),
.io_in_970(dataIn[970]),
.io_in_971(dataIn[971]),
.io_in_972(dataIn[972]),
.io_in_973(dataIn[973]),
.io_in_974(dataIn[974]),
.io_in_975(dataIn[975]),
.io_in_976(dataIn[976]),
.io_in_977(dataIn[977]),
.io_in_978(dataIn[978]),
.io_in_979(dataIn[979]),
.io_in_980(dataIn[980]),
.io_in_981(dataIn[981]),
.io_in_982(dataIn[982]),
.io_in_983(dataIn[983]),
.io_in_984(dataIn[984]),
.io_in_985(dataIn[985]),
.io_in_986(dataIn[986]),
.io_in_987(dataIn[987]),
.io_in_988(dataIn[988]),
.io_in_989(dataIn[989]),
.io_in_990(dataIn[990]),
.io_in_991(dataIn[991]),
.io_in_992(dataIn[992]),
.io_in_993(dataIn[993]),
.io_in_994(dataIn[994]),
.io_in_995(dataIn[995]),
.io_in_996(dataIn[996]),
.io_in_997(dataIn[997]),
.io_in_998(dataIn[998]),
.io_in_999(dataIn[999]),
.io_in_1000(dataIn[1000]),
.io_in_1001(dataIn[1001]),
.io_in_1002(dataIn[1002]),
.io_in_1003(dataIn[1003]),
.io_in_1004(dataIn[1004]),
.io_in_1005(dataIn[1005]),
.io_in_1006(dataIn[1006]),
.io_in_1007(dataIn[1007]),
.io_in_1008(dataIn[1008]),
.io_in_1009(dataIn[1009]),
.io_in_1010(dataIn[1010]),
.io_in_1011(dataIn[1011]),
.io_in_1012(dataIn[1012]),
.io_in_1013(dataIn[1013]),
.io_in_1014(dataIn[1014]),
.io_in_1015(dataIn[1015]),
.io_in_1016(dataIn[1016]),
.io_in_1017(dataIn[1017]),
.io_in_1018(dataIn[1018]),
.io_in_1019(dataIn[1019]),
.io_in_1020(dataIn[1020]),
.io_in_1021(dataIn[1021]),
.io_in_1022(dataIn[1022]),
.io_in_1023(dataIn[1023]),
.io_in_1024(dataIn[1024]),
.io_in_1025(dataIn[1025]),
.io_in_1026(dataIn[1026]),
.io_in_1027(dataIn[1027]),
.io_in_1028(dataIn[1028]),
.io_in_1029(dataIn[1029]),
.io_in_1030(dataIn[1030]),
.io_in_1031(dataIn[1031]),
.io_in_1032(dataIn[1032]),
.io_in_1033(dataIn[1033]),
.io_in_1034(dataIn[1034]),
.io_in_1035(dataIn[1035]),
.io_in_1036(dataIn[1036]),
.io_in_1037(dataIn[1037]),
.io_in_1038(dataIn[1038]),
.io_in_1039(dataIn[1039]),
.io_in_1040(dataIn[1040]),
.io_in_1041(dataIn[1041]),
.io_in_1042(dataIn[1042]),
.io_in_1043(dataIn[1043]),
.io_in_1044(dataIn[1044]),
.io_in_1045(dataIn[1045]),
.io_in_1046(dataIn[1046]),
.io_in_1047(dataIn[1047]),
.io_in_1048(dataIn[1048]),
.io_in_1049(dataIn[1049]),
.io_in_1050(dataIn[1050]),
.io_in_1051(dataIn[1051]),
.io_in_1052(dataIn[1052]),
.io_in_1053(dataIn[1053]),
.io_in_1054(dataIn[1054]),
.io_in_1055(dataIn[1055]),
.io_in_1056(dataIn[1056]),
.io_in_1057(dataIn[1057]),
.io_in_1058(dataIn[1058]),
.io_in_1059(dataIn[1059]),
.io_in_1060(dataIn[1060]),
.io_in_1061(dataIn[1061]),
.io_in_1062(dataIn[1062]),
.io_in_1063(dataIn[1063]),
.io_in_1064(dataIn[1064]),
.io_in_1065(dataIn[1065]),
.io_in_1066(dataIn[1066]),
.io_in_1067(dataIn[1067]),
.io_in_1068(dataIn[1068]),
.io_in_1069(dataIn[1069]),
.io_in_1070(dataIn[1070]),
.io_in_1071(dataIn[1071]),
.io_in_1072(dataIn[1072]),
.io_in_1073(dataIn[1073]),
.io_in_1074(dataIn[1074]),
.io_in_1075(dataIn[1075]),
.io_in_1076(dataIn[1076]),
.io_in_1077(dataIn[1077]),
.io_in_1078(dataIn[1078]),
.io_in_1079(dataIn[1079]),
.io_in_1080(dataIn[1080]),
.io_in_1081(dataIn[1081]),
.io_in_1082(dataIn[1082]),
.io_in_1083(dataIn[1083]),
.io_in_1084(dataIn[1084]),
.io_in_1085(dataIn[1085]),
.io_in_1086(dataIn[1086]),
.io_in_1087(dataIn[1087]),
.io_in_1088(dataIn[1088]),
.io_in_1089(dataIn[1089]),
.io_in_1090(dataIn[1090]),
.io_in_1091(dataIn[1091]),
.io_in_1092(dataIn[1092]),
.io_in_1093(dataIn[1093]),
.io_in_1094(dataIn[1094]),
.io_in_1095(dataIn[1095]),
.io_in_1096(dataIn[1096]),
.io_in_1097(dataIn[1097]),
.io_in_1098(dataIn[1098]),
.io_in_1099(dataIn[1099]),
.io_in_1100(dataIn[1100]),
.io_in_1101(dataIn[1101]),
.io_in_1102(dataIn[1102]),
.io_in_1103(dataIn[1103]),
.io_in_1104(dataIn[1104]),
.io_in_1105(dataIn[1105]),
.io_in_1106(dataIn[1106]),
.io_in_1107(dataIn[1107]),
.io_in_1108(dataIn[1108]),
.io_in_1109(dataIn[1109]),
.io_in_1110(dataIn[1110]),
.io_in_1111(dataIn[1111]),
.io_in_1112(dataIn[1112]),
.io_in_1113(dataIn[1113]),
.io_in_1114(dataIn[1114]),
.io_in_1115(dataIn[1115]),
.io_in_1116(dataIn[1116]),
.io_in_1117(dataIn[1117]),
.io_in_1118(dataIn[1118]),
.io_in_1119(dataIn[1119]),
.io_in_1120(dataIn[1120]),
.io_in_1121(dataIn[1121]),
.io_in_1122(dataIn[1122]),
.io_in_1123(dataIn[1123]),
.io_in_1124(dataIn[1124]),
.io_in_1125(dataIn[1125]),
.io_in_1126(dataIn[1126]),
.io_in_1127(dataIn[1127]),
.io_in_1128(dataIn[1128]),
.io_in_1129(dataIn[1129]),
.io_in_1130(dataIn[1130]),
.io_in_1131(dataIn[1131]),
.io_in_1132(dataIn[1132]),
.io_in_1133(dataIn[1133]),
.io_in_1134(dataIn[1134]),
.io_in_1135(dataIn[1135]),
.io_in_1136(dataIn[1136]),
.io_in_1137(dataIn[1137]),
.io_in_1138(dataIn[1138]),
.io_in_1139(dataIn[1139]),
.io_in_1140(dataIn[1140]),
.io_in_1141(dataIn[1141]),
.io_in_1142(dataIn[1142]),
.io_in_1143(dataIn[1143]),
.io_in_1144(dataIn[1144]),
.io_in_1145(dataIn[1145]),
.io_in_1146(dataIn[1146]),
.io_in_1147(dataIn[1147]),
.io_in_1148(dataIn[1148]),
.io_in_1149(dataIn[1149]),
.io_in_1150(dataIn[1150]),
.io_in_1151(dataIn[1151]),
.io_in_1152(dataIn[1152]),
.io_in_1153(dataIn[1153]),
.io_in_1154(dataIn[1154]),
.io_in_1155(dataIn[1155]),
.io_in_1156(dataIn[1156]),
.io_in_1157(dataIn[1157]),
.io_in_1158(dataIn[1158]),
.io_in_1159(dataIn[1159]),
.io_in_1160(dataIn[1160]),
.io_in_1161(dataIn[1161]),
.io_in_1162(dataIn[1162]),
.io_in_1163(dataIn[1163]),
.io_in_1164(dataIn[1164]),
.io_in_1165(dataIn[1165]),
.io_in_1166(dataIn[1166]),
.io_in_1167(dataIn[1167]),
.io_in_1168(dataIn[1168]),
.io_in_1169(dataIn[1169]),
.io_in_1170(dataIn[1170]),
.io_in_1171(dataIn[1171]),
.io_in_1172(dataIn[1172]),
.io_in_1173(dataIn[1173]),
.io_in_1174(dataIn[1174]),
.io_in_1175(dataIn[1175]),
.io_in_1176(dataIn[1176]),
.io_in_1177(dataIn[1177]),
.io_in_1178(dataIn[1178]),
.io_in_1179(dataIn[1179]),
.io_in_1180(dataIn[1180]),
.io_in_1181(dataIn[1181]),
.io_in_1182(dataIn[1182]),
.io_in_1183(dataIn[1183]),
.io_in_1184(dataIn[1184]),
.io_in_1185(dataIn[1185]),
.io_in_1186(dataIn[1186]),
.io_in_1187(dataIn[1187]),
.io_in_1188(dataIn[1188]),
.io_in_1189(dataIn[1189]),
.io_in_1190(dataIn[1190]),
.io_in_1191(dataIn[1191]),
.io_in_1192(dataIn[1192]),
.io_in_1193(dataIn[1193]),
.io_in_1194(dataIn[1194]),
.io_in_1195(dataIn[1195]),
.io_in_1196(dataIn[1196]),
.io_in_1197(dataIn[1197]),
.io_in_1198(dataIn[1198]),
.io_in_1199(dataIn[1199]),
.io_in_1200(dataIn[1200]),
.io_in_1201(dataIn[1201]),
.io_in_1202(dataIn[1202]),
.io_in_1203(dataIn[1203]),
.io_in_1204(dataIn[1204]),
.io_in_1205(dataIn[1205]),
.io_in_1206(dataIn[1206]),
.io_in_1207(dataIn[1207]),
.io_in_1208(dataIn[1208]),
.io_in_1209(dataIn[1209]),
.io_in_1210(dataIn[1210]),
.io_in_1211(dataIn[1211]),
.io_in_1212(dataIn[1212]),
.io_in_1213(dataIn[1213]),
.io_in_1214(dataIn[1214]),
.io_in_1215(dataIn[1215]),
.io_in_1216(dataIn[1216]),
.io_in_1217(dataIn[1217]),
.io_in_1218(dataIn[1218]),
.io_in_1219(dataIn[1219]),
.io_in_1220(dataIn[1220]),
.io_in_1221(dataIn[1221]),
.io_in_1222(dataIn[1222]),
.io_in_1223(dataIn[1223]),
.io_in_1224(dataIn[1224]),
.io_in_1225(dataIn[1225]),
.io_in_1226(dataIn[1226]),
.io_in_1227(dataIn[1227]),
.io_in_1228(dataIn[1228]),
.io_in_1229(dataIn[1229]),
.io_in_1230(dataIn[1230]),
.io_in_1231(dataIn[1231]),
.io_in_1232(dataIn[1232]),
.io_in_1233(dataIn[1233]),
.io_in_1234(dataIn[1234]),
.io_in_1235(dataIn[1235]),
.io_in_1236(dataIn[1236]),
.io_in_1237(dataIn[1237]),
.io_in_1238(dataIn[1238]),
.io_in_1239(dataIn[1239]),
.io_in_1240(dataIn[1240]),
.io_in_1241(dataIn[1241]),
.io_in_1242(dataIn[1242]),
.io_in_1243(dataIn[1243]),
.io_in_1244(dataIn[1244]),
.io_in_1245(dataIn[1245]),
.io_in_1246(dataIn[1246]),
.io_in_1247(dataIn[1247]),
.io_in_1248(dataIn[1248]),
.io_in_1249(dataIn[1249]),
.io_in_1250(dataIn[1250]),
.io_in_1251(dataIn[1251]),
.io_in_1252(dataIn[1252]),
.io_in_1253(dataIn[1253]),
.io_in_1254(dataIn[1254]),
.io_in_1255(dataIn[1255]),
.io_in_1256(dataIn[1256]),
.io_in_1257(dataIn[1257]),
.io_in_1258(dataIn[1258]),
.io_in_1259(dataIn[1259]),
.io_in_1260(dataIn[1260]),
.io_in_1261(dataIn[1261]),
.io_in_1262(dataIn[1262]),
.io_in_1263(dataIn[1263]),
.io_in_1264(dataIn[1264]),
.io_in_1265(dataIn[1265]),
.io_in_1266(dataIn[1266]),
.io_in_1267(dataIn[1267]),
.io_in_1268(dataIn[1268]),
.io_in_1269(dataIn[1269]),
.io_in_1270(dataIn[1270]),
.io_in_1271(dataIn[1271]),
.io_in_1272(dataIn[1272]),
.io_in_1273(dataIn[1273]),
.io_in_1274(dataIn[1274]),
.io_in_1275(dataIn[1275]),
.io_in_1276(dataIn[1276]),
.io_in_1277(dataIn[1277]),
.io_in_1278(dataIn[1278]),
.io_in_1279(dataIn[1279]),
.io_in_1280(dataIn[1280]),
.io_in_1281(dataIn[1281]),
.io_in_1282(dataIn[1282]),
.io_in_1283(dataIn[1283]),
.io_in_1284(dataIn[1284]),
.io_in_1285(dataIn[1285]),
.io_in_1286(dataIn[1286]),
.io_in_1287(dataIn[1287]),
.io_in_1288(dataIn[1288]),
.io_in_1289(dataIn[1289]),
.io_in_1290(dataIn[1290]),
.io_in_1291(dataIn[1291]),
.io_in_1292(dataIn[1292]),
.io_in_1293(dataIn[1293]),
.io_in_1294(dataIn[1294]),
.io_in_1295(dataIn[1295]),
.io_in_1296(dataIn[1296]),
.io_in_1297(dataIn[1297]),
.io_in_1298(dataIn[1298]),
.io_in_1299(dataIn[1299]),
.io_in_1300(dataIn[1300]),
.io_in_1301(dataIn[1301]),
.io_in_1302(dataIn[1302]),
.io_in_1303(dataIn[1303]),
.io_in_1304(dataIn[1304]),
.io_in_1305(dataIn[1305]),
.io_in_1306(dataIn[1306]),
.io_in_1307(dataIn[1307]),
.io_in_1308(dataIn[1308]),
.io_in_1309(dataIn[1309]),
.io_in_1310(dataIn[1310]),
.io_in_1311(dataIn[1311]),
.io_in_1312(dataIn[1312]),
.io_in_1313(dataIn[1313]),
.io_in_1314(dataIn[1314]),
.io_in_1315(dataIn[1315]),
.io_in_1316(dataIn[1316]),
.io_in_1317(dataIn[1317]),
.io_in_1318(dataIn[1318]),
.io_in_1319(dataIn[1319]),
.io_in_1320(dataIn[1320]),
.io_in_1321(dataIn[1321]),
.io_in_1322(dataIn[1322]),
.io_in_1323(dataIn[1323]),
.io_in_1324(dataIn[1324]),
.io_in_1325(dataIn[1325]),
.io_in_1326(dataIn[1326]),
.io_in_1327(dataIn[1327]),
.io_in_1328(dataIn[1328]),
.io_in_1329(dataIn[1329]),
.io_in_1330(dataIn[1330]),
.io_in_1331(dataIn[1331]),
.io_in_1332(dataIn[1332]),
.io_in_1333(dataIn[1333]),
.io_in_1334(dataIn[1334]),
.io_in_1335(dataIn[1335]),
.io_in_1336(dataIn[1336]),
.io_in_1337(dataIn[1337]),
.io_in_1338(dataIn[1338]),
.io_in_1339(dataIn[1339]),
.io_in_1340(dataIn[1340]),
.io_in_1341(dataIn[1341]),
.io_in_1342(dataIn[1342]),
.io_in_1343(dataIn[1343]),
.io_in_1344(dataIn[1344]),
.io_in_1345(dataIn[1345]),
.io_in_1346(dataIn[1346]),
.io_in_1347(dataIn[1347]),
.io_in_1348(dataIn[1348]),
.io_in_1349(dataIn[1349]),
.io_in_1350(dataIn[1350]),
.io_in_1351(dataIn[1351]),
.io_in_1352(dataIn[1352]),
.io_in_1353(dataIn[1353]),
.io_in_1354(dataIn[1354]),
.io_in_1355(dataIn[1355]),
.io_in_1356(dataIn[1356]),
.io_in_1357(dataIn[1357]),
.io_in_1358(dataIn[1358]),
.io_in_1359(dataIn[1359]),
.io_in_1360(dataIn[1360]),
.io_in_1361(dataIn[1361]),
.io_in_1362(dataIn[1362]),
.io_in_1363(dataIn[1363]),
.io_in_1364(dataIn[1364]),
.io_in_1365(dataIn[1365]),
.io_in_1366(dataIn[1366]),
.io_in_1367(dataIn[1367]),
.io_in_1368(dataIn[1368]),
.io_in_1369(dataIn[1369]),
.io_in_1370(dataIn[1370]),
.io_in_1371(dataIn[1371]),
.io_in_1372(dataIn[1372]),
.io_in_1373(dataIn[1373]),
.io_in_1374(dataIn[1374]),
.io_in_1375(dataIn[1375]),
.io_in_1376(dataIn[1376]),
.io_in_1377(dataIn[1377]),
.io_in_1378(dataIn[1378]),
.io_in_1379(dataIn[1379]),
.io_in_1380(dataIn[1380]),
.io_in_1381(dataIn[1381]),
.io_in_1382(dataIn[1382]),
.io_in_1383(dataIn[1383]),
.io_in_1384(dataIn[1384]),
.io_in_1385(dataIn[1385]),
.io_in_1386(dataIn[1386]),
.io_in_1387(dataIn[1387]),
.io_in_1388(dataIn[1388]),
.io_in_1389(dataIn[1389]),
.io_in_1390(dataIn[1390]),
.io_in_1391(dataIn[1391]),
.io_in_1392(dataIn[1392]),
.io_in_1393(dataIn[1393]),
.io_in_1394(dataIn[1394]),
.io_in_1395(dataIn[1395]),
.io_in_1396(dataIn[1396]),
.io_in_1397(dataIn[1397]),
.io_in_1398(dataIn[1398]),
.io_in_1399(dataIn[1399]),
.io_in_1400(dataIn[1400]),
.io_in_1401(dataIn[1401]),
.io_in_1402(dataIn[1402]),
.io_in_1403(dataIn[1403]),
.io_in_1404(dataIn[1404]),
.io_in_1405(dataIn[1405]),
.io_in_1406(dataIn[1406]),
.io_in_1407(dataIn[1407]),
.io_in_1408(dataIn[1408]),
.io_in_1409(dataIn[1409]),
.io_in_1410(dataIn[1410]),
.io_in_1411(dataIn[1411]),
.io_in_1412(dataIn[1412]),
.io_in_1413(dataIn[1413]),
.io_in_1414(dataIn[1414]),
.io_in_1415(dataIn[1415]),
.io_in_1416(dataIn[1416]),
.io_in_1417(dataIn[1417]),
.io_in_1418(dataIn[1418]),
.io_in_1419(dataIn[1419]),
.io_in_1420(dataIn[1420]),
.io_in_1421(dataIn[1421]),
.io_in_1422(dataIn[1422]),
.io_in_1423(dataIn[1423]),
.io_in_1424(dataIn[1424]),
.io_in_1425(dataIn[1425]),
.io_in_1426(dataIn[1426]),
.io_in_1427(dataIn[1427]),
.io_in_1428(dataIn[1428]),
.io_in_1429(dataIn[1429]),
.io_in_1430(dataIn[1430]),
.io_in_1431(dataIn[1431]),
.io_in_1432(dataIn[1432]),
.io_in_1433(dataIn[1433]),
.io_in_1434(dataIn[1434]),
.io_in_1435(dataIn[1435]),
.io_in_1436(dataIn[1436]),
.io_in_1437(dataIn[1437]),
.io_in_1438(dataIn[1438]),
.io_in_1439(dataIn[1439]),
.io_in_1440(dataIn[1440]),
.io_in_1441(dataIn[1441]),
.io_in_1442(dataIn[1442]),
.io_in_1443(dataIn[1443]),
.io_in_1444(dataIn[1444]),
.io_in_1445(dataIn[1445]),
.io_in_1446(dataIn[1446]),
.io_in_1447(dataIn[1447]),
.io_in_1448(dataIn[1448]),
.io_in_1449(dataIn[1449]),
.io_in_1450(dataIn[1450]),
.io_in_1451(dataIn[1451]),
.io_in_1452(dataIn[1452]),
.io_in_1453(dataIn[1453]),
.io_in_1454(dataIn[1454]),
.io_in_1455(dataIn[1455]),
.io_in_1456(dataIn[1456]),
.io_in_1457(dataIn[1457]),
.io_in_1458(dataIn[1458]),
.io_in_1459(dataIn[1459]),
.io_in_1460(dataIn[1460]),
.io_in_1461(dataIn[1461]),
.io_in_1462(dataIn[1462]),
.io_in_1463(dataIn[1463]),
.io_in_1464(dataIn[1464]),
.io_in_1465(dataIn[1465]),
.io_in_1466(dataIn[1466]),
.io_in_1467(dataIn[1467]),
.io_in_1468(dataIn[1468]),
.io_in_1469(dataIn[1469]),
.io_in_1470(dataIn[1470]),
.io_in_1471(dataIn[1471]),
.io_in_1472(dataIn[1472]),
.io_in_1473(dataIn[1473]),
.io_in_1474(dataIn[1474]),
.io_in_1475(dataIn[1475]),
.io_in_1476(dataIn[1476]),
.io_in_1477(dataIn[1477]),
.io_in_1478(dataIn[1478]),
.io_in_1479(dataIn[1479]),
.io_in_1480(dataIn[1480]),
.io_in_1481(dataIn[1481]),
.io_in_1482(dataIn[1482]),
.io_in_1483(dataIn[1483]),
.io_in_1484(dataIn[1484]),
.io_in_1485(dataIn[1485]),
.io_in_1486(dataIn[1486]),
.io_in_1487(dataIn[1487]),
.io_in_1488(dataIn[1488]),
.io_in_1489(dataIn[1489]),
.io_in_1490(dataIn[1490]),
.io_in_1491(dataIn[1491]),
.io_in_1492(dataIn[1492]),
.io_in_1493(dataIn[1493]),
.io_in_1494(dataIn[1494]),
.io_in_1495(dataIn[1495]),
.io_in_1496(dataIn[1496]),
.io_in_1497(dataIn[1497]),
.io_in_1498(dataIn[1498]),
.io_in_1499(dataIn[1499]),
.io_in_1500(dataIn[1500]),
.io_in_1501(dataIn[1501]),
.io_in_1502(dataIn[1502]),
.io_in_1503(dataIn[1503]),
.io_in_1504(dataIn[1504]),
.io_in_1505(dataIn[1505]),
.io_in_1506(dataIn[1506]),
.io_in_1507(dataIn[1507]),
.io_in_1508(dataIn[1508]),
.io_in_1509(dataIn[1509]),
.io_in_1510(dataIn[1510]),
.io_in_1511(dataIn[1511]),
.io_in_1512(dataIn[1512]),
.io_in_1513(dataIn[1513]),
.io_in_1514(dataIn[1514]),
.io_in_1515(dataIn[1515]),
.io_in_1516(dataIn[1516]),
.io_in_1517(dataIn[1517]),
.io_in_1518(dataIn[1518]),
.io_in_1519(dataIn[1519]),
.io_in_1520(dataIn[1520]),
.io_in_1521(dataIn[1521]),
.io_in_1522(dataIn[1522]),
.io_in_1523(dataIn[1523]),
.io_in_1524(dataIn[1524]),
.io_in_1525(dataIn[1525]),
.io_in_1526(dataIn[1526]),
.io_in_1527(dataIn[1527]),
.io_in_1528(dataIn[1528]),
.io_in_1529(dataIn[1529]),
.io_in_1530(dataIn[1530]),
.io_in_1531(dataIn[1531]),
.io_in_1532(dataIn[1532]),
.io_in_1533(dataIn[1533]),
.io_in_1534(dataIn[1534]),
.io_in_1535(dataIn[1535]),
.io_in_1536(dataIn[1536]),
.io_in_1537(dataIn[1537]),
.io_in_1538(dataIn[1538]),
.io_in_1539(dataIn[1539]),
.io_in_1540(dataIn[1540]),
.io_in_1541(dataIn[1541]),
.io_in_1542(dataIn[1542]),
.io_in_1543(dataIn[1543]),
.io_in_1544(dataIn[1544]),
.io_in_1545(dataIn[1545]),
.io_in_1546(dataIn[1546]),
.io_in_1547(dataIn[1547]),
.io_in_1548(dataIn[1548]),
.io_in_1549(dataIn[1549]),
.io_in_1550(dataIn[1550]),
.io_in_1551(dataIn[1551]),
.io_in_1552(dataIn[1552]),
.io_in_1553(dataIn[1553]),
.io_in_1554(dataIn[1554]),
.io_in_1555(dataIn[1555]),
.io_in_1556(dataIn[1556]),
.io_in_1557(dataIn[1557]),
.io_in_1558(dataIn[1558]),
.io_in_1559(dataIn[1559]),
.io_in_1560(dataIn[1560]),
.io_in_1561(dataIn[1561]),
.io_in_1562(dataIn[1562]),
.io_in_1563(dataIn[1563]),
.io_in_1564(dataIn[1564]),
.io_in_1565(dataIn[1565]),
.io_in_1566(dataIn[1566]),
.io_in_1567(dataIn[1567]),
.io_in_1568(dataIn[1568]),
.io_in_1569(dataIn[1569]),
.io_in_1570(dataIn[1570]),
.io_in_1571(dataIn[1571]),
.io_in_1572(dataIn[1572]),
.io_in_1573(dataIn[1573]),
.io_in_1574(dataIn[1574]),
.io_in_1575(dataIn[1575]),
.io_in_1576(dataIn[1576]),
.io_in_1577(dataIn[1577]),
.io_in_1578(dataIn[1578]),
.io_in_1579(dataIn[1579]),
.io_in_1580(dataIn[1580]),
.io_in_1581(dataIn[1581]),
.io_in_1582(dataIn[1582]),
.io_in_1583(dataIn[1583]),
.io_in_1584(dataIn[1584]),
.io_in_1585(dataIn[1585]),
.io_in_1586(dataIn[1586]),
.io_in_1587(dataIn[1587]),
.io_in_1588(dataIn[1588]),
.io_in_1589(dataIn[1589]),
.io_in_1590(dataIn[1590]),
.io_in_1591(dataIn[1591]),
.io_in_1592(dataIn[1592]),
.io_in_1593(dataIn[1593]),
.io_in_1594(dataIn[1594]),
.io_in_1595(dataIn[1595]),
.io_in_1596(dataIn[1596]),
.io_in_1597(dataIn[1597]),
.io_in_1598(dataIn[1598]),
.io_in_1599(dataIn[1599]),
.io_in_1600(dataIn[1600]),
.io_in_1601(dataIn[1601]),
.io_in_1602(dataIn[1602]),
.io_in_1603(dataIn[1603]),
.io_in_1604(dataIn[1604]),
.io_in_1605(dataIn[1605]),
.io_in_1606(dataIn[1606]),
.io_in_1607(dataIn[1607]),
.io_in_1608(dataIn[1608]),
.io_in_1609(dataIn[1609]),
.io_in_1610(dataIn[1610]),
.io_in_1611(dataIn[1611]),
.io_in_1612(dataIn[1612]),
.io_in_1613(dataIn[1613]),
.io_in_1614(dataIn[1614]),
.io_in_1615(dataIn[1615]),
.io_in_1616(dataIn[1616]),
.io_in_1617(dataIn[1617]),
.io_in_1618(dataIn[1618]),
.io_in_1619(dataIn[1619]),
.io_in_1620(dataIn[1620]),
.io_in_1621(dataIn[1621]),
.io_in_1622(dataIn[1622]),
.io_in_1623(dataIn[1623]),
.io_in_1624(dataIn[1624]),
.io_in_1625(dataIn[1625]),
.io_in_1626(dataIn[1626]),
.io_in_1627(dataIn[1627]),
.io_in_1628(dataIn[1628]),
.io_in_1629(dataIn[1629]),
.io_in_1630(dataIn[1630]),
.io_in_1631(dataIn[1631]),
.io_in_1632(dataIn[1632]),
.io_in_1633(dataIn[1633]),
.io_in_1634(dataIn[1634]),
.io_in_1635(dataIn[1635]),
.io_in_1636(dataIn[1636]),
.io_in_1637(dataIn[1637]),
.io_in_1638(dataIn[1638]),
.io_in_1639(dataIn[1639]),
.io_in_1640(dataIn[1640]),
.io_in_1641(dataIn[1641]),
.io_in_1642(dataIn[1642]),
.io_in_1643(dataIn[1643]),
.io_in_1644(dataIn[1644]),
.io_in_1645(dataIn[1645]),
.io_in_1646(dataIn[1646]),
.io_in_1647(dataIn[1647]),
.io_in_1648(dataIn[1648]),
.io_in_1649(dataIn[1649]),
.io_in_1650(dataIn[1650]),
.io_in_1651(dataIn[1651]),
.io_in_1652(dataIn[1652]),
.io_in_1653(dataIn[1653]),
.io_in_1654(dataIn[1654]),
.io_in_1655(dataIn[1655]),
.io_in_1656(dataIn[1656]),
.io_in_1657(dataIn[1657]),
.io_in_1658(dataIn[1658]),
.io_in_1659(dataIn[1659]),
.io_in_1660(dataIn[1660]),
.io_in_1661(dataIn[1661]),
.io_in_1662(dataIn[1662]),
.io_in_1663(dataIn[1663]),
.io_in_1664(dataIn[1664]),
.io_in_1665(dataIn[1665]),
.io_in_1666(dataIn[1666]),
.io_in_1667(dataIn[1667]),
.io_in_1668(dataIn[1668]),
.io_in_1669(dataIn[1669]),
.io_in_1670(dataIn[1670]),
.io_in_1671(dataIn[1671]),
.io_in_1672(dataIn[1672]),
.io_in_1673(dataIn[1673]),
.io_in_1674(dataIn[1674]),
.io_in_1675(dataIn[1675]),
.io_in_1676(dataIn[1676]),
.io_in_1677(dataIn[1677]),
.io_in_1678(dataIn[1678]),
.io_in_1679(dataIn[1679]),
.io_in_1680(dataIn[1680]),
.io_in_1681(dataIn[1681]),
.io_in_1682(dataIn[1682]),
.io_in_1683(dataIn[1683]),
.io_in_1684(dataIn[1684]),
.io_in_1685(dataIn[1685]),
.io_in_1686(dataIn[1686]),
.io_in_1687(dataIn[1687]),
.io_in_1688(dataIn[1688]),
.io_in_1689(dataIn[1689]),
.io_in_1690(dataIn[1690]),
.io_in_1691(dataIn[1691]),
.io_in_1692(dataIn[1692]),
.io_in_1693(dataIn[1693]),
.io_in_1694(dataIn[1694]),
.io_in_1695(dataIn[1695]),
.io_in_1696(dataIn[1696]),
.io_in_1697(dataIn[1697]),
.io_in_1698(dataIn[1698]),
.io_in_1699(dataIn[1699]),
.io_in_1700(dataIn[1700]),
.io_in_1701(dataIn[1701]),
.io_in_1702(dataIn[1702]),
.io_in_1703(dataIn[1703]),
.io_in_1704(dataIn[1704]),
.io_in_1705(dataIn[1705]),
.io_in_1706(dataIn[1706]),
.io_in_1707(dataIn[1707]),
.io_in_1708(dataIn[1708]),
.io_in_1709(dataIn[1709]),
.io_in_1710(dataIn[1710]),
.io_in_1711(dataIn[1711]),
.io_in_1712(dataIn[1712]),
.io_in_1713(dataIn[1713]),
.io_in_1714(dataIn[1714]),
.io_in_1715(dataIn[1715]),
.io_in_1716(dataIn[1716]),
.io_in_1717(dataIn[1717]),
.io_in_1718(dataIn[1718]),
.io_in_1719(dataIn[1719]),
.io_in_1720(dataIn[1720]),
.io_in_1721(dataIn[1721]),
.io_in_1722(dataIn[1722]),
.io_in_1723(dataIn[1723]),
.io_in_1724(dataIn[1724]),
.io_in_1725(dataIn[1725]),
.io_in_1726(dataIn[1726]),
.io_in_1727(dataIn[1727]),
.io_in_1728(dataIn[1728]),
.io_in_1729(dataIn[1729]),
.io_in_1730(dataIn[1730]),
.io_in_1731(dataIn[1731]),
.io_in_1732(dataIn[1732]),
.io_in_1733(dataIn[1733]),
.io_in_1734(dataIn[1734]),
.io_in_1735(dataIn[1735]),
.io_in_1736(dataIn[1736]),
.io_in_1737(dataIn[1737]),
.io_in_1738(dataIn[1738]),
.io_in_1739(dataIn[1739]),
.io_in_1740(dataIn[1740]),
.io_in_1741(dataIn[1741]),
.io_in_1742(dataIn[1742]),
.io_in_1743(dataIn[1743]),
.io_in_1744(dataIn[1744]),
.io_in_1745(dataIn[1745]),
.io_in_1746(dataIn[1746]),
.io_in_1747(dataIn[1747]),
.io_in_1748(dataIn[1748]),
.io_in_1749(dataIn[1749]),
.io_in_1750(dataIn[1750]),
.io_in_1751(dataIn[1751]),
.io_in_1752(dataIn[1752]),
.io_in_1753(dataIn[1753]),
.io_in_1754(dataIn[1754]),
.io_in_1755(dataIn[1755]),
.io_in_1756(dataIn[1756]),
.io_in_1757(dataIn[1757]),
.io_in_1758(dataIn[1758]),
.io_in_1759(dataIn[1759]),
.io_in_1760(dataIn[1760]),
.io_in_1761(dataIn[1761]),
.io_in_1762(dataIn[1762]),
.io_in_1763(dataIn[1763]),
.io_in_1764(dataIn[1764]),
.io_in_1765(dataIn[1765]),
.io_in_1766(dataIn[1766]),
.io_in_1767(dataIn[1767]),
.io_in_1768(dataIn[1768]),
.io_in_1769(dataIn[1769]),
.io_in_1770(dataIn[1770]),
.io_in_1771(dataIn[1771]),
.io_in_1772(dataIn[1772]),
.io_in_1773(dataIn[1773]),
.io_in_1774(dataIn[1774]),
.io_in_1775(dataIn[1775]),
.io_in_1776(dataIn[1776]),
.io_in_1777(dataIn[1777]),
.io_in_1778(dataIn[1778]),
.io_in_1779(dataIn[1779]),
.io_in_1780(dataIn[1780]),
.io_in_1781(dataIn[1781]),
.io_in_1782(dataIn[1782]),
.io_in_1783(dataIn[1783]),
.io_in_1784(dataIn[1784]),
.io_in_1785(dataIn[1785]),
.io_in_1786(dataIn[1786]),
.io_in_1787(dataIn[1787]),
.io_in_1788(dataIn[1788]),
.io_in_1789(dataIn[1789]),
.io_in_1790(dataIn[1790]),
.io_in_1791(dataIn[1791]),
.io_in_1792(dataIn[1792]),
.io_in_1793(dataIn[1793]),
.io_in_1794(dataIn[1794]),
.io_in_1795(dataIn[1795]),
.io_in_1796(dataIn[1796]),
.io_in_1797(dataIn[1797]),
.io_in_1798(dataIn[1798]),
.io_in_1799(dataIn[1799]),
.io_in_1800(dataIn[1800]),
.io_in_1801(dataIn[1801]),
.io_in_1802(dataIn[1802]),
.io_in_1803(dataIn[1803]),
.io_in_1804(dataIn[1804]),
.io_in_1805(dataIn[1805]),
.io_in_1806(dataIn[1806]),
.io_in_1807(dataIn[1807]),
.io_in_1808(dataIn[1808]),
.io_in_1809(dataIn[1809]),
.io_in_1810(dataIn[1810]),
.io_in_1811(dataIn[1811]),
.io_in_1812(dataIn[1812]),
.io_in_1813(dataIn[1813]),
.io_in_1814(dataIn[1814]),
.io_in_1815(dataIn[1815]),
.io_in_1816(dataIn[1816]),
.io_in_1817(dataIn[1817]),
.io_in_1818(dataIn[1818]),
.io_in_1819(dataIn[1819]),
.io_in_1820(dataIn[1820]),
.io_in_1821(dataIn[1821]),
.io_in_1822(dataIn[1822]),
.io_in_1823(dataIn[1823]),
.io_in_1824(dataIn[1824]),
.io_in_1825(dataIn[1825]),
.io_in_1826(dataIn[1826]),
.io_in_1827(dataIn[1827]),
.io_in_1828(dataIn[1828]),
.io_in_1829(dataIn[1829]),
.io_in_1830(dataIn[1830]),
.io_in_1831(dataIn[1831]),
.io_in_1832(dataIn[1832]),
.io_in_1833(dataIn[1833]),
.io_in_1834(dataIn[1834]),
.io_in_1835(dataIn[1835]),
.io_in_1836(dataIn[1836]),
.io_in_1837(dataIn[1837]),
.io_in_1838(dataIn[1838]),
.io_in_1839(dataIn[1839]),
.io_in_1840(dataIn[1840]),
.io_in_1841(dataIn[1841]),
.io_in_1842(dataIn[1842]),
.io_in_1843(dataIn[1843]),
.io_in_1844(dataIn[1844]),
.io_in_1845(dataIn[1845]),
.io_in_1846(dataIn[1846]),
.io_in_1847(dataIn[1847]),
.io_in_1848(dataIn[1848]),
.io_in_1849(dataIn[1849]),
.io_in_1850(dataIn[1850]),
.io_in_1851(dataIn[1851]),
.io_in_1852(dataIn[1852]),
.io_in_1853(dataIn[1853]),
.io_in_1854(dataIn[1854]),
.io_in_1855(dataIn[1855]),
.io_in_1856(dataIn[1856]),
.io_in_1857(dataIn[1857]),
.io_in_1858(dataIn[1858]),
.io_in_1859(dataIn[1859]),
.io_in_1860(dataIn[1860]),
.io_in_1861(dataIn[1861]),
.io_in_1862(dataIn[1862]),
.io_in_1863(dataIn[1863]),
.io_in_1864(dataIn[1864]),
.io_in_1865(dataIn[1865]),
.io_in_1866(dataIn[1866]),
.io_in_1867(dataIn[1867]),
.io_in_1868(dataIn[1868]),
.io_in_1869(dataIn[1869]),
.io_in_1870(dataIn[1870]),
.io_in_1871(dataIn[1871]),
.io_in_1872(dataIn[1872]),
.io_in_1873(dataIn[1873]),
.io_in_1874(dataIn[1874]),
.io_in_1875(dataIn[1875]),
.io_in_1876(dataIn[1876]),
.io_in_1877(dataIn[1877]),
.io_in_1878(dataIn[1878]),
.io_in_1879(dataIn[1879]),
.io_in_1880(dataIn[1880]),
.io_in_1881(dataIn[1881]),
.io_in_1882(dataIn[1882]),
.io_in_1883(dataIn[1883]),
.io_in_1884(dataIn[1884]),
.io_in_1885(dataIn[1885]),
.io_in_1886(dataIn[1886]),
.io_in_1887(dataIn[1887]),
.io_in_1888(dataIn[1888]),
.io_in_1889(dataIn[1889]),
.io_in_1890(dataIn[1890]),
.io_in_1891(dataIn[1891]),
.io_in_1892(dataIn[1892]),
.io_in_1893(dataIn[1893]),
.io_in_1894(dataIn[1894]),
.io_in_1895(dataIn[1895]),
.io_in_1896(dataIn[1896]),
.io_in_1897(dataIn[1897]),
.io_in_1898(dataIn[1898]),
.io_in_1899(dataIn[1899]),
.io_in_1900(dataIn[1900]),
.io_in_1901(dataIn[1901]),
.io_in_1902(dataIn[1902]),
.io_in_1903(dataIn[1903]),
.io_in_1904(dataIn[1904]),
.io_in_1905(dataIn[1905]),
.io_in_1906(dataIn[1906]),
.io_in_1907(dataIn[1907]),
.io_in_1908(dataIn[1908]),
.io_in_1909(dataIn[1909]),
.io_in_1910(dataIn[1910]),
.io_in_1911(dataIn[1911]),
.io_in_1912(dataIn[1912]),
.io_in_1913(dataIn[1913]),
.io_in_1914(dataIn[1914]),
.io_in_1915(dataIn[1915]),
.io_in_1916(dataIn[1916]),
.io_in_1917(dataIn[1917]),
.io_in_1918(dataIn[1918]),
.io_in_1919(dataIn[1919]),
.io_in_1920(dataIn[1920]),
.io_in_1921(dataIn[1921]),
.io_in_1922(dataIn[1922]),
.io_in_1923(dataIn[1923]),
.io_in_1924(dataIn[1924]),
.io_in_1925(dataIn[1925]),
.io_in_1926(dataIn[1926]),
.io_in_1927(dataIn[1927]),
.io_in_1928(dataIn[1928]),
.io_in_1929(dataIn[1929]),
.io_in_1930(dataIn[1930]),
.io_in_1931(dataIn[1931]),
.io_in_1932(dataIn[1932]),
.io_in_1933(dataIn[1933]),
.io_in_1934(dataIn[1934]),
.io_in_1935(dataIn[1935]),
.io_in_1936(dataIn[1936]),
.io_in_1937(dataIn[1937]),
.io_in_1938(dataIn[1938]),
.io_in_1939(dataIn[1939]),
.io_in_1940(dataIn[1940]),
.io_in_1941(dataIn[1941]),
.io_in_1942(dataIn[1942]),
.io_in_1943(dataIn[1943]),
.io_in_1944(dataIn[1944]),
.io_in_1945(dataIn[1945]),
.io_in_1946(dataIn[1946]),
.io_in_1947(dataIn[1947]),
.io_in_1948(dataIn[1948]),
.io_in_1949(dataIn[1949]),
.io_in_1950(dataIn[1950]),
.io_in_1951(dataIn[1951]),
.io_in_1952(dataIn[1952]),
.io_in_1953(dataIn[1953]),
.io_in_1954(dataIn[1954]),
.io_in_1955(dataIn[1955]),
.io_in_1956(dataIn[1956]),
.io_in_1957(dataIn[1957]),
.io_in_1958(dataIn[1958]),
.io_in_1959(dataIn[1959]),
.io_in_1960(dataIn[1960]),
.io_in_1961(dataIn[1961]),
.io_in_1962(dataIn[1962]),
.io_in_1963(dataIn[1963]),
.io_in_1964(dataIn[1964]),
.io_in_1965(dataIn[1965]),
.io_in_1966(dataIn[1966]),
.io_in_1967(dataIn[1967]),
.io_in_1968(dataIn[1968]),
.io_in_1969(dataIn[1969]),
.io_in_1970(dataIn[1970]),
.io_in_1971(dataIn[1971]),
.io_in_1972(dataIn[1972]),
.io_in_1973(dataIn[1973]),
.io_in_1974(dataIn[1974]),
.io_in_1975(dataIn[1975]),
.io_in_1976(dataIn[1976]),
.io_in_1977(dataIn[1977]),
.io_in_1978(dataIn[1978]),
.io_in_1979(dataIn[1979]),
.io_in_1980(dataIn[1980]),
.io_in_1981(dataIn[1981]),
.io_in_1982(dataIn[1982]),
.io_in_1983(dataIn[1983]),
.io_in_1984(dataIn[1984]),
.io_in_1985(dataIn[1985]),
.io_in_1986(dataIn[1986]),
.io_in_1987(dataIn[1987]),
.io_in_1988(dataIn[1988]),
.io_in_1989(dataIn[1989]),
.io_in_1990(dataIn[1990]),
.io_in_1991(dataIn[1991]),
.io_in_1992(dataIn[1992]),
.io_in_1993(dataIn[1993]),
.io_in_1994(dataIn[1994]),
.io_in_1995(dataIn[1995]),
.io_in_1996(dataIn[1996]),
.io_in_1997(dataIn[1997]),
.io_in_1998(dataIn[1998]),
.io_in_1999(dataIn[1999]),
.io_in_2000(dataIn[2000]),
.io_in_2001(dataIn[2001]),
.io_in_2002(dataIn[2002]),
.io_in_2003(dataIn[2003]),
.io_in_2004(dataIn[2004]),
.io_in_2005(dataIn[2005]),
.io_in_2006(dataIn[2006]),
.io_in_2007(dataIn[2007]),
.io_in_2008(dataIn[2008]),
.io_in_2009(dataIn[2009]),
.io_in_2010(dataIn[2010]),
.io_in_2011(dataIn[2011]),
.io_in_2012(dataIn[2012]),
.io_in_2013(dataIn[2013]),
.io_in_2014(dataIn[2014]),
.io_in_2015(dataIn[2015]),
.io_in_2016(dataIn[2016]),
.io_in_2017(dataIn[2017]),
.io_in_2018(dataIn[2018]),
.io_in_2019(dataIn[2019]),
.io_in_2020(dataIn[2020]),
.io_in_2021(dataIn[2021]),
.io_in_2022(dataIn[2022]),
.io_in_2023(dataIn[2023]),
.io_in_2024(dataIn[2024]),
.io_in_2025(dataIn[2025]),
.io_in_2026(dataIn[2026]),
.io_in_2027(dataIn[2027]),
.io_in_2028(dataIn[2028]),
.io_in_2029(dataIn[2029]),
.io_in_2030(dataIn[2030]),
.io_in_2031(dataIn[2031]),
.io_in_2032(dataIn[2032]),
.io_in_2033(dataIn[2033]),
.io_in_2034(dataIn[2034]),
.io_in_2035(dataIn[2035]),
.io_in_2036(dataIn[2036]),
.io_in_2037(dataIn[2037]),
.io_in_2038(dataIn[2038]),
.io_in_2039(dataIn[2039]),
.io_in_2040(dataIn[2040]),
.io_in_2041(dataIn[2041]),
.io_in_2042(dataIn[2042]),
.io_in_2043(dataIn[2043]),
.io_in_2044(dataIn[2044]),
.io_in_2045(dataIn[2045]),
.io_in_2046(dataIn[2046]),
.io_in_2047(dataIn[2047]),
.io_in_2048(dataIn[2048]),
.io_in_2049(dataIn[2049]),
.io_in_2050(dataIn[2050]),
.io_in_2051(dataIn[2051]),
.io_in_2052(dataIn[2052]),
.io_in_2053(dataIn[2053]),
.io_in_2054(dataIn[2054]),
.io_in_2055(dataIn[2055]),
.io_in_2056(dataIn[2056]),
.io_in_2057(dataIn[2057]),
.io_in_2058(dataIn[2058]),
.io_in_2059(dataIn[2059]),
.io_in_2060(dataIn[2060]),
.io_in_2061(dataIn[2061]),
.io_in_2062(dataIn[2062]),
.io_in_2063(dataIn[2063]),
.io_in_2064(dataIn[2064]),
.io_in_2065(dataIn[2065]),
.io_in_2066(dataIn[2066]),
.io_in_2067(dataIn[2067]),
.io_in_2068(dataIn[2068]),
.io_in_2069(dataIn[2069]),
.io_in_2070(dataIn[2070]),
.io_in_2071(dataIn[2071]),
.io_in_2072(dataIn[2072]),
.io_in_2073(dataIn[2073]),
.io_in_2074(dataIn[2074]),
.io_in_2075(dataIn[2075]),
.io_in_2076(dataIn[2076]),
.io_in_2077(dataIn[2077]),
.io_in_2078(dataIn[2078]),
.io_in_2079(dataIn[2079]),
.io_in_2080(dataIn[2080]),
.io_in_2081(dataIn[2081]),
.io_in_2082(dataIn[2082]),
.io_in_2083(dataIn[2083]),
.io_in_2084(dataIn[2084]),
.io_in_2085(dataIn[2085]),
.io_in_2086(dataIn[2086]),
.io_in_2087(dataIn[2087]),
.io_in_2088(dataIn[2088]),
.io_in_2089(dataIn[2089]),
.io_in_2090(dataIn[2090]),
.io_in_2091(dataIn[2091]),
.io_in_2092(dataIn[2092]),
.io_in_2093(dataIn[2093]),
.io_in_2094(dataIn[2094]),
.io_in_2095(dataIn[2095]),
.io_in_2096(dataIn[2096]),
.io_in_2097(dataIn[2097]),
.io_in_2098(dataIn[2098]),
.io_in_2099(dataIn[2099]),
.io_in_2100(dataIn[2100]),
.io_in_2101(dataIn[2101]),
.io_in_2102(dataIn[2102]),
.io_in_2103(dataIn[2103]),
.io_in_2104(dataIn[2104]),
.io_in_2105(dataIn[2105]),
.io_in_2106(dataIn[2106]),
.io_in_2107(dataIn[2107]),
.io_in_2108(dataIn[2108]),
.io_in_2109(dataIn[2109]),
.io_in_2110(dataIn[2110]),
.io_in_2111(dataIn[2111]),
.io_in_2112(dataIn[2112]),
.io_in_2113(dataIn[2113]),
.io_in_2114(dataIn[2114]),
.io_in_2115(dataIn[2115]),
.io_in_2116(dataIn[2116]),
.io_in_2117(dataIn[2117]),
.io_in_2118(dataIn[2118]),
.io_in_2119(dataIn[2119]),
.io_in_2120(dataIn[2120]),
.io_in_2121(dataIn[2121]),
.io_in_2122(dataIn[2122]),
.io_in_2123(dataIn[2123]),
.io_in_2124(dataIn[2124]),
.io_in_2125(dataIn[2125]),
.io_in_2126(dataIn[2126]),
.io_in_2127(dataIn[2127]),
.io_in_2128(dataIn[2128]),
.io_in_2129(dataIn[2129]),
.io_in_2130(dataIn[2130]),
.io_in_2131(dataIn[2131]),
.io_in_2132(dataIn[2132]),
.io_in_2133(dataIn[2133]),
.io_in_2134(dataIn[2134]),
.io_in_2135(dataIn[2135]),
.io_in_2136(dataIn[2136]),
.io_in_2137(dataIn[2137]),
.io_in_2138(dataIn[2138]),
.io_in_2139(dataIn[2139]),
.io_in_2140(dataIn[2140]),
.io_in_2141(dataIn[2141]),
.io_in_2142(dataIn[2142]),
.io_in_2143(dataIn[2143]),
.io_in_2144(dataIn[2144]),
.io_in_2145(dataIn[2145]),
.io_in_2146(dataIn[2146]),
.io_in_2147(dataIn[2147]),
.io_in_2148(dataIn[2148]),
.io_in_2149(dataIn[2149]),
.io_in_2150(dataIn[2150]),
.io_in_2151(dataIn[2151]),
.io_in_2152(dataIn[2152]),
.io_in_2153(dataIn[2153]),
.io_in_2154(dataIn[2154]),
.io_in_2155(dataIn[2155]),
.io_in_2156(dataIn[2156]),
.io_in_2157(dataIn[2157]),
.io_in_2158(dataIn[2158]),
.io_in_2159(dataIn[2159]),
.io_in_2160(dataIn[2160]),
.io_in_2161(dataIn[2161]),
.io_in_2162(dataIn[2162]),
.io_in_2163(dataIn[2163]),
.io_in_2164(dataIn[2164]),
.io_in_2165(dataIn[2165]),
.io_in_2166(dataIn[2166]),
.io_in_2167(dataIn[2167]),
.io_in_2168(dataIn[2168]),
.io_in_2169(dataIn[2169]),
.io_in_2170(dataIn[2170]),
.io_in_2171(dataIn[2171]),
.io_in_2172(dataIn[2172]),
.io_in_2173(dataIn[2173]),
.io_in_2174(dataIn[2174]),
.io_in_2175(dataIn[2175]),
.io_in_2176(dataIn[2176]),
.io_in_2177(dataIn[2177]),
.io_in_2178(dataIn[2178]),
.io_in_2179(dataIn[2179]),
.io_in_2180(dataIn[2180]),
.io_in_2181(dataIn[2181]),
.io_in_2182(dataIn[2182]),
.io_in_2183(dataIn[2183]),
.io_in_2184(dataIn[2184]),
.io_in_2185(dataIn[2185]),
.io_in_2186(dataIn[2186]),
.io_in_2187(dataIn[2187]),
.io_in_2188(dataIn[2188]),
.io_in_2189(dataIn[2189]),
.io_in_2190(dataIn[2190]),
.io_in_2191(dataIn[2191]),
.io_in_2192(dataIn[2192]),
.io_in_2193(dataIn[2193]),
.io_in_2194(dataIn[2194]),
.io_in_2195(dataIn[2195]),
.io_in_2196(dataIn[2196]),
.io_in_2197(dataIn[2197]),
.io_in_2198(dataIn[2198]),
.io_in_2199(dataIn[2199]),
.io_in_2200(dataIn[2200]),
.io_in_2201(dataIn[2201]),
.io_in_2202(dataIn[2202]),
.io_in_2203(dataIn[2203]),
.io_in_2204(dataIn[2204]),
.io_in_2205(dataIn[2205]),
.io_in_2206(dataIn[2206]),
.io_in_2207(dataIn[2207]),
.io_in_2208(dataIn[2208]),
.io_in_2209(dataIn[2209]),
.io_in_2210(dataIn[2210]),
.io_in_2211(dataIn[2211]),
.io_in_2212(dataIn[2212]),
.io_in_2213(dataIn[2213]),
.io_in_2214(dataIn[2214]),
.io_in_2215(dataIn[2215]),
.io_in_2216(dataIn[2216]),
.io_in_2217(dataIn[2217]),
.io_in_2218(dataIn[2218]),
.io_in_2219(dataIn[2219]),
.io_in_2220(dataIn[2220]),
.io_in_2221(dataIn[2221]),
.io_in_2222(dataIn[2222]),
.io_in_2223(dataIn[2223]),
.io_in_2224(dataIn[2224]),
.io_in_2225(dataIn[2225]),
.io_in_2226(dataIn[2226]),
.io_in_2227(dataIn[2227]),
.io_in_2228(dataIn[2228]),
.io_in_2229(dataIn[2229]),
.io_in_2230(dataIn[2230]),
.io_in_2231(dataIn[2231]),
.io_in_2232(dataIn[2232]),
.io_in_2233(dataIn[2233]),
.io_in_2234(dataIn[2234]),
.io_in_2235(dataIn[2235]),
.io_in_2236(dataIn[2236]),
.io_in_2237(dataIn[2237]),
.io_in_2238(dataIn[2238]),
.io_in_2239(dataIn[2239]),
.io_in_2240(dataIn[2240]),
.io_in_2241(dataIn[2241]),
.io_in_2242(dataIn[2242]),
.io_in_2243(dataIn[2243]),
.io_in_2244(dataIn[2244]),
.io_in_2245(dataIn[2245]),
.io_in_2246(dataIn[2246]),
.io_in_2247(dataIn[2247]),
.io_in_2248(dataIn[2248]),
.io_in_2249(dataIn[2249]),
.io_in_2250(dataIn[2250]),
.io_in_2251(dataIn[2251]),
.io_in_2252(dataIn[2252]),
.io_in_2253(dataIn[2253]),
.io_in_2254(dataIn[2254]),
.io_in_2255(dataIn[2255]),
.io_in_2256(dataIn[2256]),
.io_in_2257(dataIn[2257]),
.io_in_2258(dataIn[2258]),
.io_in_2259(dataIn[2259]),
.io_in_2260(dataIn[2260]),
.io_in_2261(dataIn[2261]),
.io_in_2262(dataIn[2262]),
.io_in_2263(dataIn[2263]),
.io_in_2264(dataIn[2264]),
.io_in_2265(dataIn[2265]),
.io_in_2266(dataIn[2266]),
.io_in_2267(dataIn[2267]),
.io_in_2268(dataIn[2268]),
.io_in_2269(dataIn[2269]),
.io_in_2270(dataIn[2270]),
.io_in_2271(dataIn[2271]),
.io_in_2272(dataIn[2272]),
.io_in_2273(dataIn[2273]),
.io_in_2274(dataIn[2274]),
.io_in_2275(dataIn[2275]),
.io_in_2276(dataIn[2276]),
.io_in_2277(dataIn[2277]),
.io_in_2278(dataIn[2278]),
.io_in_2279(dataIn[2279]),
.io_in_2280(dataIn[2280]),
.io_in_2281(dataIn[2281]),
.io_in_2282(dataIn[2282]),
.io_in_2283(dataIn[2283]),
.io_in_2284(dataIn[2284]),
.io_in_2285(dataIn[2285]),
.io_in_2286(dataIn[2286]),
.io_in_2287(dataIn[2287]),
.io_in_2288(dataIn[2288]),
.io_in_2289(dataIn[2289]),
.io_in_2290(dataIn[2290]),
.io_in_2291(dataIn[2291]),
.io_in_2292(dataIn[2292]),
.io_in_2293(dataIn[2293]),
.io_in_2294(dataIn[2294]),
.io_in_2295(dataIn[2295]),
.io_in_2296(dataIn[2296]),
.io_in_2297(dataIn[2297]),
.io_in_2298(dataIn[2298]),
.io_in_2299(dataIn[2299]),
.io_in_2300(dataIn[2300]),
.io_in_2301(dataIn[2301]),
.io_in_2302(dataIn[2302]),
.io_in_2303(dataIn[2303]),
.io_in_2304(dataIn[2304]),
.io_in_2305(dataIn[2305]),
.io_in_2306(dataIn[2306]),
.io_in_2307(dataIn[2307]),
.io_in_2308(dataIn[2308]),
.io_in_2309(dataIn[2309]),
.io_in_2310(dataIn[2310]),
.io_in_2311(dataIn[2311]),
.io_in_2312(dataIn[2312]),
.io_in_2313(dataIn[2313]),
.io_in_2314(dataIn[2314]),
.io_in_2315(dataIn[2315]),
.io_in_2316(dataIn[2316]),
.io_in_2317(dataIn[2317]),
.io_in_2318(dataIn[2318]),
.io_in_2319(dataIn[2319]),
.io_in_2320(dataIn[2320]),
.io_in_2321(dataIn[2321]),
.io_in_2322(dataIn[2322]),
.io_in_2323(dataIn[2323]),
.io_in_2324(dataIn[2324]),
.io_in_2325(dataIn[2325]),
.io_in_2326(dataIn[2326]),
.io_in_2327(dataIn[2327]),
.io_in_2328(dataIn[2328]),
.io_in_2329(dataIn[2329]),
.io_in_2330(dataIn[2330]),
.io_in_2331(dataIn[2331]),
.io_in_2332(dataIn[2332]),
.io_in_2333(dataIn[2333]),
.io_in_2334(dataIn[2334]),
.io_in_2335(dataIn[2335]),
.io_in_2336(dataIn[2336]),
.io_in_2337(dataIn[2337]),
.io_in_2338(dataIn[2338]),
.io_in_2339(dataIn[2339]),
.io_in_2340(dataIn[2340]),
.io_in_2341(dataIn[2341]),
.io_in_2342(dataIn[2342]),
.io_in_2343(dataIn[2343]),
.io_in_2344(dataIn[2344]),
.io_in_2345(dataIn[2345]),
.io_in_2346(dataIn[2346]),
.io_in_2347(dataIn[2347]),
.io_in_2348(dataIn[2348]),
.io_in_2349(dataIn[2349]),
.io_in_2350(dataIn[2350]),
.io_in_2351(dataIn[2351]),
.io_in_2352(dataIn[2352]),
.io_in_2353(dataIn[2353]),
.io_in_2354(dataIn[2354]),
.io_in_2355(dataIn[2355]),
.io_in_2356(dataIn[2356]),
.io_in_2357(dataIn[2357]),
.io_in_2358(dataIn[2358]),
.io_in_2359(dataIn[2359]),
.io_in_2360(dataIn[2360]),
.io_in_2361(dataIn[2361]),
.io_in_2362(dataIn[2362]),
.io_in_2363(dataIn[2363]),
.io_in_2364(dataIn[2364]),
.io_in_2365(dataIn[2365]),
.io_in_2366(dataIn[2366]),
.io_in_2367(dataIn[2367]),
.io_in_2368(dataIn[2368]),
.io_in_2369(dataIn[2369]),
.io_in_2370(dataIn[2370]),
.io_in_2371(dataIn[2371]),
.io_in_2372(dataIn[2372]),
.io_in_2373(dataIn[2373]),
.io_in_2374(dataIn[2374]),
.io_in_2375(dataIn[2375]),
.io_in_2376(dataIn[2376]),
.io_in_2377(dataIn[2377]),
.io_in_2378(dataIn[2378]),
.io_in_2379(dataIn[2379]),
.io_in_2380(dataIn[2380]),
.io_in_2381(dataIn[2381]),
.io_in_2382(dataIn[2382]),
.io_in_2383(dataIn[2383]),
.io_in_2384(dataIn[2384]),
.io_in_2385(dataIn[2385]),
.io_in_2386(dataIn[2386]),
.io_in_2387(dataIn[2387]),
.io_in_2388(dataIn[2388]),
.io_in_2389(dataIn[2389]),
.io_in_2390(dataIn[2390]),
.io_in_2391(dataIn[2391]),
.io_in_2392(dataIn[2392]),
.io_in_2393(dataIn[2393]),
.io_in_2394(dataIn[2394]),
.io_in_2395(dataIn[2395]),
.io_in_2396(dataIn[2396]),
.io_in_2397(dataIn[2397]),
.io_in_2398(dataIn[2398]),
.io_in_2399(dataIn[2399]),
.io_in_2400(dataIn[2400]),
.io_in_2401(dataIn[2401]),
.io_in_2402(dataIn[2402]),
.io_in_2403(dataIn[2403]),
.io_in_2404(dataIn[2404]),
.io_in_2405(dataIn[2405]),
.io_in_2406(dataIn[2406]),
.io_in_2407(dataIn[2407]),
.io_in_2408(dataIn[2408]),
.io_in_2409(dataIn[2409]),
.io_in_2410(dataIn[2410]),
.io_in_2411(dataIn[2411]),
.io_in_2412(dataIn[2412]),
.io_in_2413(dataIn[2413]),
.io_in_2414(dataIn[2414]),
.io_in_2415(dataIn[2415]),
.io_in_2416(dataIn[2416]),
.io_in_2417(dataIn[2417]),
.io_in_2418(dataIn[2418]),
.io_in_2419(dataIn[2419]),
.io_in_2420(dataIn[2420]),
.io_in_2421(dataIn[2421]),
.io_in_2422(dataIn[2422]),
.io_in_2423(dataIn[2423]),
.io_in_2424(dataIn[2424]),
.io_in_2425(dataIn[2425]),
.io_in_2426(dataIn[2426]),
.io_in_2427(dataIn[2427]),
.io_in_2428(dataIn[2428]),
.io_in_2429(dataIn[2429]),
.io_in_2430(dataIn[2430]),
.io_in_2431(dataIn[2431]),
.io_in_2432(dataIn[2432]),
.io_in_2433(dataIn[2433]),
.io_in_2434(dataIn[2434]),
.io_in_2435(dataIn[2435]),
.io_in_2436(dataIn[2436]),
.io_in_2437(dataIn[2437]),
.io_in_2438(dataIn[2438]),
.io_in_2439(dataIn[2439]),
.io_in_2440(dataIn[2440]),
.io_in_2441(dataIn[2441]),
.io_in_2442(dataIn[2442]),
.io_in_2443(dataIn[2443]),
.io_in_2444(dataIn[2444]),
.io_in_2445(dataIn[2445]),
.io_in_2446(dataIn[2446]),
.io_in_2447(dataIn[2447]),
.io_in_2448(dataIn[2448]),
.io_in_2449(dataIn[2449]),
.io_in_2450(dataIn[2450]),
.io_in_2451(dataIn[2451]),
.io_in_2452(dataIn[2452]),
.io_in_2453(dataIn[2453]),
.io_in_2454(dataIn[2454]),
.io_in_2455(dataIn[2455]),
.io_in_2456(dataIn[2456]),
.io_in_2457(dataIn[2457]),
.io_in_2458(dataIn[2458]),
.io_in_2459(dataIn[2459]),
.io_in_2460(dataIn[2460]),
.io_in_2461(dataIn[2461]),
.io_in_2462(dataIn[2462]),
.io_in_2463(dataIn[2463]),
.io_in_2464(dataIn[2464]),
.io_in_2465(dataIn[2465]),
.io_in_2466(dataIn[2466]),
.io_in_2467(dataIn[2467]),
.io_in_2468(dataIn[2468]),
.io_in_2469(dataIn[2469]),
.io_in_2470(dataIn[2470]),
.io_in_2471(dataIn[2471]),
.io_in_2472(dataIn[2472]),
.io_in_2473(dataIn[2473]),
.io_in_2474(dataIn[2474]),
.io_in_2475(dataIn[2475]),
.io_in_2476(dataIn[2476]),
.io_in_2477(dataIn[2477]),
.io_in_2478(dataIn[2478]),
.io_in_2479(dataIn[2479]),
.io_in_2480(dataIn[2480]),
.io_in_2481(dataIn[2481]),
.io_in_2482(dataIn[2482]),
.io_in_2483(dataIn[2483]),
.io_in_2484(dataIn[2484]),
.io_in_2485(dataIn[2485]),
.io_in_2486(dataIn[2486]),
.io_in_2487(dataIn[2487]),
.io_in_2488(dataIn[2488]),
.io_in_2489(dataIn[2489]),
.io_in_2490(dataIn[2490]),
.io_in_2491(dataIn[2491]),
.io_in_2492(dataIn[2492]),
.io_in_2493(dataIn[2493]),
.io_in_2494(dataIn[2494]),
.io_in_2495(dataIn[2495]),
.io_in_2496(dataIn[2496]),
.io_in_2497(dataIn[2497]),
.io_in_2498(dataIn[2498]),
.io_in_2499(dataIn[2499]),
.io_in_2500(dataIn[2500]),
.io_in_2501(dataIn[2501]),
.io_in_2502(dataIn[2502]),
.io_in_2503(dataIn[2503]),
.io_in_2504(dataIn[2504]),
.io_in_2505(dataIn[2505]),
.io_in_2506(dataIn[2506]),
.io_in_2507(dataIn[2507]),
.io_in_2508(dataIn[2508]),
.io_in_2509(dataIn[2509]),
.io_in_2510(dataIn[2510]),
.io_in_2511(dataIn[2511]),
.io_in_2512(dataIn[2512]),
.io_in_2513(dataIn[2513]),
.io_in_2514(dataIn[2514]),
.io_in_2515(dataIn[2515]),
.io_in_2516(dataIn[2516]),
.io_in_2517(dataIn[2517]),
.io_in_2518(dataIn[2518]),
.io_in_2519(dataIn[2519]),
.io_in_2520(dataIn[2520]),
.io_in_2521(dataIn[2521]),
.io_in_2522(dataIn[2522]),
.io_in_2523(dataIn[2523]),
.io_in_2524(dataIn[2524]),
.io_in_2525(dataIn[2525]),
.io_in_2526(dataIn[2526]),
.io_in_2527(dataIn[2527]),
.io_in_2528(dataIn[2528]),
.io_in_2529(dataIn[2529]),
.io_in_2530(dataIn[2530]),
.io_in_2531(dataIn[2531]),
.io_in_2532(dataIn[2532]),
.io_in_2533(dataIn[2533]),
.io_in_2534(dataIn[2534]),
.io_in_2535(dataIn[2535]),
.io_in_2536(dataIn[2536]),
.io_in_2537(dataIn[2537]),
.io_in_2538(dataIn[2538]),
.io_in_2539(dataIn[2539]),
.io_in_2540(dataIn[2540]),
.io_in_2541(dataIn[2541]),
.io_in_2542(dataIn[2542]),
.io_in_2543(dataIn[2543]),
.io_in_2544(dataIn[2544]),
.io_in_2545(dataIn[2545]),
.io_in_2546(dataIn[2546]),
.io_in_2547(dataIn[2547]),
.io_in_2548(dataIn[2548]),
.io_in_2549(dataIn[2549]),
.io_in_2550(dataIn[2550]),
.io_in_2551(dataIn[2551]),
.io_in_2552(dataIn[2552]),
.io_in_2553(dataIn[2553]),
.io_in_2554(dataIn[2554]),
.io_in_2555(dataIn[2555]),
.io_in_2556(dataIn[2556]),
.io_in_2557(dataIn[2557]),
.io_in_2558(dataIn[2558]),
.io_in_2559(dataIn[2559]),
.io_in_2560(dataIn[2560]),
.io_in_2561(dataIn[2561]),
.io_in_2562(dataIn[2562]),
.io_in_2563(dataIn[2563]),
.io_in_2564(dataIn[2564]),
.io_in_2565(dataIn[2565]),
.io_in_2566(dataIn[2566]),
.io_in_2567(dataIn[2567]),
.io_in_2568(dataIn[2568]),
.io_in_2569(dataIn[2569]),
.io_in_2570(dataIn[2570]),
.io_in_2571(dataIn[2571]),
.io_in_2572(dataIn[2572]),
.io_in_2573(dataIn[2573]),
.io_in_2574(dataIn[2574]),
.io_in_2575(dataIn[2575]),
.io_in_2576(dataIn[2576]),
.io_in_2577(dataIn[2577]),
.io_in_2578(dataIn[2578]),
.io_in_2579(dataIn[2579]),
.io_in_2580(dataIn[2580]),
.io_in_2581(dataIn[2581]),
.io_in_2582(dataIn[2582]),
.io_in_2583(dataIn[2583]),
.io_in_2584(dataIn[2584]),
.io_in_2585(dataIn[2585]),
.io_in_2586(dataIn[2586]),
.io_in_2587(dataIn[2587]),
.io_in_2588(dataIn[2588]),
.io_in_2589(dataIn[2589]),
.io_in_2590(dataIn[2590]),
.io_in_2591(dataIn[2591]),
.io_in_2592(dataIn[2592]),
.io_in_2593(dataIn[2593]),
.io_in_2594(dataIn[2594]),
.io_in_2595(dataIn[2595]),
.io_in_2596(dataIn[2596]),
.io_in_2597(dataIn[2597]),
.io_in_2598(dataIn[2598]),
.io_in_2599(dataIn[2599]),
.io_in_2600(dataIn[2600]),
.io_in_2601(dataIn[2601]),
.io_in_2602(dataIn[2602]),
.io_in_2603(dataIn[2603]),
.io_in_2604(dataIn[2604]),
.io_in_2605(dataIn[2605]),
.io_in_2606(dataIn[2606]),
.io_in_2607(dataIn[2607]),
.io_in_2608(dataIn[2608]),
.io_in_2609(dataIn[2609]),
.io_in_2610(dataIn[2610]),
.io_in_2611(dataIn[2611]),
.io_in_2612(dataIn[2612]),
.io_in_2613(dataIn[2613]),
.io_in_2614(dataIn[2614]),
.io_in_2615(dataIn[2615]),
.io_in_2616(dataIn[2616]),
.io_in_2617(dataIn[2617]),
.io_in_2618(dataIn[2618]),
.io_in_2619(dataIn[2619]),
.io_in_2620(dataIn[2620]),
.io_in_2621(dataIn[2621]),
.io_in_2622(dataIn[2622]),
.io_in_2623(dataIn[2623]),
.io_in_2624(dataIn[2624]),
.io_in_2625(dataIn[2625]),
.io_in_2626(dataIn[2626]),
.io_in_2627(dataIn[2627]),
.io_in_2628(dataIn[2628]),
.io_in_2629(dataIn[2629]),
.io_in_2630(dataIn[2630]),
.io_in_2631(dataIn[2631]),
.io_in_2632(dataIn[2632]),
.io_in_2633(dataIn[2633]),
.io_in_2634(dataIn[2634]),
.io_in_2635(dataIn[2635]),
.io_in_2636(dataIn[2636]),
.io_in_2637(dataIn[2637]),
.io_in_2638(dataIn[2638]),
.io_in_2639(dataIn[2639]),
.io_in_2640(dataIn[2640]),
.io_in_2641(dataIn[2641]),
.io_in_2642(dataIn[2642]),
.io_in_2643(dataIn[2643]),
.io_in_2644(dataIn[2644]),
.io_in_2645(dataIn[2645]),
.io_in_2646(dataIn[2646]),
.io_in_2647(dataIn[2647]),
.io_in_2648(dataIn[2648]),
.io_in_2649(dataIn[2649]),
.io_in_2650(dataIn[2650]),
.io_in_2651(dataIn[2651]),
.io_in_2652(dataIn[2652]),
.io_in_2653(dataIn[2653]),
.io_in_2654(dataIn[2654]),
.io_in_2655(dataIn[2655]),
.io_in_2656(dataIn[2656]),
.io_in_2657(dataIn[2657]),
.io_in_2658(dataIn[2658]),
.io_in_2659(dataIn[2659]),
.io_in_2660(dataIn[2660]),
.io_in_2661(dataIn[2661]),
.io_in_2662(dataIn[2662]),
.io_in_2663(dataIn[2663]),
.io_in_2664(dataIn[2664]),
.io_in_2665(dataIn[2665]),
.io_in_2666(dataIn[2666]),
.io_in_2667(dataIn[2667]),
.io_in_2668(dataIn[2668]),
.io_in_2669(dataIn[2669]),
.io_in_2670(dataIn[2670]),
.io_in_2671(dataIn[2671]),
.io_in_2672(dataIn[2672]),
.io_in_2673(dataIn[2673]),
.io_in_2674(dataIn[2674]),
.io_in_2675(dataIn[2675]),
.io_in_2676(dataIn[2676]),
.io_in_2677(dataIn[2677]),
.io_in_2678(dataIn[2678]),
.io_in_2679(dataIn[2679]),
.io_in_2680(dataIn[2680]),
.io_in_2681(dataIn[2681]),
.io_in_2682(dataIn[2682]),
.io_in_2683(dataIn[2683]),
.io_in_2684(dataIn[2684]),
.io_in_2685(dataIn[2685]),
.io_in_2686(dataIn[2686]),
.io_in_2687(dataIn[2687]),
.io_in_2688(dataIn[2688]),
.io_in_2689(dataIn[2689]),
.io_in_2690(dataIn[2690]),
.io_in_2691(dataIn[2691]),
.io_in_2692(dataIn[2692]),
.io_in_2693(dataIn[2693]),
.io_in_2694(dataIn[2694]),
.io_in_2695(dataIn[2695]),
.io_in_2696(dataIn[2696]),
.io_in_2697(dataIn[2697]),
.io_in_2698(dataIn[2698]),
.io_in_2699(dataIn[2699]),
.io_in_2700(dataIn[2700]),
.io_in_2701(dataIn[2701]),
.io_in_2702(dataIn[2702]),
.io_in_2703(dataIn[2703]),
.io_in_2704(dataIn[2704]),
.io_in_2705(dataIn[2705]),
.io_in_2706(dataIn[2706]),
.io_in_2707(dataIn[2707]),
.io_in_2708(dataIn[2708]),
.io_in_2709(dataIn[2709]),
.io_in_2710(dataIn[2710]),
.io_in_2711(dataIn[2711]),
.io_in_2712(dataIn[2712]),
.io_in_2713(dataIn[2713]),
.io_in_2714(dataIn[2714]),
.io_in_2715(dataIn[2715]),
.io_in_2716(dataIn[2716]),
.io_in_2717(dataIn[2717]),
.io_in_2718(dataIn[2718]),
.io_in_2719(dataIn[2719]),
.io_in_2720(dataIn[2720]),
.io_in_2721(dataIn[2721]),
.io_in_2722(dataIn[2722]),
.io_in_2723(dataIn[2723]),
.io_in_2724(dataIn[2724]),
.io_in_2725(dataIn[2725]),
.io_in_2726(dataIn[2726]),
.io_in_2727(dataIn[2727]),
.io_in_2728(dataIn[2728]),
.io_in_2729(dataIn[2729]),
.io_in_2730(dataIn[2730]),
.io_in_2731(dataIn[2731]),
.io_in_2732(dataIn[2732]),
.io_in_2733(dataIn[2733]),
.io_in_2734(dataIn[2734]),
.io_in_2735(dataIn[2735]),
.io_in_2736(dataIn[2736]),
.io_in_2737(dataIn[2737]),
.io_in_2738(dataIn[2738]),
.io_in_2739(dataIn[2739]),
.io_in_2740(dataIn[2740]),
.io_in_2741(dataIn[2741]),
.io_in_2742(dataIn[2742]),
.io_in_2743(dataIn[2743]),
.io_in_2744(dataIn[2744]),
.io_in_2745(dataIn[2745]),
.io_in_2746(dataIn[2746]),
.io_in_2747(dataIn[2747]),
.io_in_2748(dataIn[2748]),
.io_in_2749(dataIn[2749]),
.io_in_2750(dataIn[2750]),
.io_in_2751(dataIn[2751]),
.io_in_2752(dataIn[2752]),
.io_in_2753(dataIn[2753]),
.io_in_2754(dataIn[2754]),
.io_in_2755(dataIn[2755]),
.io_in_2756(dataIn[2756]),
.io_in_2757(dataIn[2757]),
.io_in_2758(dataIn[2758]),
.io_in_2759(dataIn[2759]),
.io_in_2760(dataIn[2760]),
.io_in_2761(dataIn[2761]),
.io_in_2762(dataIn[2762]),
.io_in_2763(dataIn[2763]),
.io_in_2764(dataIn[2764]),
.io_in_2765(dataIn[2765]),
.io_in_2766(dataIn[2766]),
.io_in_2767(dataIn[2767]),
.io_in_2768(dataIn[2768]),
.io_in_2769(dataIn[2769]),
.io_in_2770(dataIn[2770]),
.io_in_2771(dataIn[2771]),
.io_in_2772(dataIn[2772]),
.io_in_2773(dataIn[2773]),
.io_in_2774(dataIn[2774]),
.io_in_2775(dataIn[2775]),
.io_in_2776(dataIn[2776]),
.io_in_2777(dataIn[2777]),
.io_in_2778(dataIn[2778]),
.io_in_2779(dataIn[2779]),
.io_in_2780(dataIn[2780]),
.io_in_2781(dataIn[2781]),
.io_in_2782(dataIn[2782]),
.io_in_2783(dataIn[2783]),
.io_in_2784(dataIn[2784]),
.io_in_2785(dataIn[2785]),
.io_in_2786(dataIn[2786]),
.io_in_2787(dataIn[2787]),
.io_in_2788(dataIn[2788]),
.io_in_2789(dataIn[2789]),
.io_in_2790(dataIn[2790]),
.io_in_2791(dataIn[2791]),
.io_in_2792(dataIn[2792]),
.io_in_2793(dataIn[2793]),
.io_in_2794(dataIn[2794]),
.io_in_2795(dataIn[2795]),
.io_in_2796(dataIn[2796]),
.io_in_2797(dataIn[2797]),
.io_in_2798(dataIn[2798]),
.io_in_2799(dataIn[2799]),
.io_in_2800(dataIn[2800]),
.io_in_2801(dataIn[2801]),
.io_in_2802(dataIn[2802]),
.io_in_2803(dataIn[2803]),
.io_in_2804(dataIn[2804]),
.io_in_2805(dataIn[2805]),
.io_in_2806(dataIn[2806]),
.io_in_2807(dataIn[2807]),
.io_in_2808(dataIn[2808]),
.io_in_2809(dataIn[2809]),
.io_in_2810(dataIn[2810]),
.io_in_2811(dataIn[2811]),
.io_in_2812(dataIn[2812]),
.io_in_2813(dataIn[2813]),
.io_in_2814(dataIn[2814]),
.io_in_2815(dataIn[2815]),
.io_in_2816(dataIn[2816]),
.io_in_2817(dataIn[2817]),
.io_in_2818(dataIn[2818]),
.io_in_2819(dataIn[2819]),
.io_in_2820(dataIn[2820]),
.io_in_2821(dataIn[2821]),
.io_in_2822(dataIn[2822]),
.io_in_2823(dataIn[2823]),
.io_in_2824(dataIn[2824]),
.io_in_2825(dataIn[2825]),
.io_in_2826(dataIn[2826]),
.io_in_2827(dataIn[2827]),
.io_in_2828(dataIn[2828]),
.io_in_2829(dataIn[2829]),
.io_in_2830(dataIn[2830]),
.io_in_2831(dataIn[2831]),
.io_in_2832(dataIn[2832]),
.io_in_2833(dataIn[2833]),
.io_in_2834(dataIn[2834]),
.io_in_2835(dataIn[2835]),
.io_in_2836(dataIn[2836]),
.io_in_2837(dataIn[2837]),
.io_in_2838(dataIn[2838]),
.io_in_2839(dataIn[2839]),
.io_in_2840(dataIn[2840]),
.io_in_2841(dataIn[2841]),
.io_in_2842(dataIn[2842]),
.io_in_2843(dataIn[2843]),
.io_in_2844(dataIn[2844]),
.io_in_2845(dataIn[2845]),
.io_in_2846(dataIn[2846]),
.io_in_2847(dataIn[2847]),
.io_in_2848(dataIn[2848]),
.io_in_2849(dataIn[2849]),
.io_in_2850(dataIn[2850]),
.io_in_2851(dataIn[2851]),
.io_in_2852(dataIn[2852]),
.io_in_2853(dataIn[2853]),
.io_in_2854(dataIn[2854]),
.io_in_2855(dataIn[2855]),
.io_in_2856(dataIn[2856]),
.io_in_2857(dataIn[2857]),
.io_in_2858(dataIn[2858]),
.io_in_2859(dataIn[2859]),
.io_in_2860(dataIn[2860]),
.io_in_2861(dataIn[2861]),
.io_in_2862(dataIn[2862]),
.io_in_2863(dataIn[2863]),
.io_in_2864(dataIn[2864]),
.io_in_2865(dataIn[2865]),
.io_in_2866(dataIn[2866]),
.io_in_2867(dataIn[2867]),
.io_in_2868(dataIn[2868]),
.io_in_2869(dataIn[2869]),
.io_in_2870(dataIn[2870]),
.io_in_2871(dataIn[2871]),
.io_in_2872(dataIn[2872]),
.io_in_2873(dataIn[2873]),
.io_in_2874(dataIn[2874]),
.io_in_2875(dataIn[2875]),
.io_in_2876(dataIn[2876]),
.io_in_2877(dataIn[2877]),
.io_in_2878(dataIn[2878]),
.io_in_2879(dataIn[2879]),
.io_in_2880(dataIn[2880]),
.io_in_2881(dataIn[2881]),
.io_in_2882(dataIn[2882]),
.io_in_2883(dataIn[2883]),
.io_in_2884(dataIn[2884]),
.io_in_2885(dataIn[2885]),
.io_in_2886(dataIn[2886]),
.io_in_2887(dataIn[2887]),
.io_in_2888(dataIn[2888]),
.io_in_2889(dataIn[2889]),
.io_in_2890(dataIn[2890]),
.io_in_2891(dataIn[2891]),
.io_in_2892(dataIn[2892]),
.io_in_2893(dataIn[2893]),
.io_in_2894(dataIn[2894]),
.io_in_2895(dataIn[2895]),
.io_in_2896(dataIn[2896]),
.io_in_2897(dataIn[2897]),
.io_in_2898(dataIn[2898]),
.io_in_2899(dataIn[2899]),
.io_in_2900(dataIn[2900]),
.io_in_2901(dataIn[2901]),
.io_in_2902(dataIn[2902]),
.io_in_2903(dataIn[2903]),
.io_in_2904(dataIn[2904]),
.io_in_2905(dataIn[2905]),
.io_in_2906(dataIn[2906]),
.io_in_2907(dataIn[2907]),
.io_in_2908(dataIn[2908]),
.io_in_2909(dataIn[2909]),
.io_in_2910(dataIn[2910]),
.io_in_2911(dataIn[2911]),
.io_in_2912(dataIn[2912]),
.io_in_2913(dataIn[2913]),
.io_in_2914(dataIn[2914]),
.io_in_2915(dataIn[2915]),
.io_in_2916(dataIn[2916]),
.io_in_2917(dataIn[2917]),
.io_in_2918(dataIn[2918]),
.io_in_2919(dataIn[2919]),
.io_in_2920(dataIn[2920]),
.io_in_2921(dataIn[2921]),
.io_in_2922(dataIn[2922]),
.io_in_2923(dataIn[2923]),
.io_in_2924(dataIn[2924]),
.io_in_2925(dataIn[2925]),
.io_in_2926(dataIn[2926]),
.io_in_2927(dataIn[2927]),
.io_in_2928(dataIn[2928]),
.io_in_2929(dataIn[2929]),
.io_in_2930(dataIn[2930]),
.io_in_2931(dataIn[2931]),
.io_in_2932(dataIn[2932]),
.io_in_2933(dataIn[2933]),
.io_in_2934(dataIn[2934]),
.io_in_2935(dataIn[2935]),
.io_in_2936(dataIn[2936]),
.io_in_2937(dataIn[2937]),
.io_in_2938(dataIn[2938]),
.io_in_2939(dataIn[2939]),
.io_in_2940(dataIn[2940]),
.io_in_2941(dataIn[2941]),
.io_in_2942(dataIn[2942]),
.io_in_2943(dataIn[2943]),
.io_in_2944(dataIn[2944]),
.io_in_2945(dataIn[2945]),
.io_in_2946(dataIn[2946]),
.io_in_2947(dataIn[2947]),
.io_in_2948(dataIn[2948]),
.io_in_2949(dataIn[2949]),
.io_in_2950(dataIn[2950]),
.io_in_2951(dataIn[2951]),
.io_in_2952(dataIn[2952]),
.io_in_2953(dataIn[2953]),
.io_in_2954(dataIn[2954]),
.io_in_2955(dataIn[2955]),
.io_in_2956(dataIn[2956]),
.io_in_2957(dataIn[2957]),
.io_in_2958(dataIn[2958]),
.io_in_2959(dataIn[2959]),
.io_in_2960(dataIn[2960]),
.io_in_2961(dataIn[2961]),
.io_in_2962(dataIn[2962]),
.io_in_2963(dataIn[2963]),
.io_in_2964(dataIn[2964]),
.io_in_2965(dataIn[2965]),
.io_in_2966(dataIn[2966]),
.io_in_2967(dataIn[2967]),
.io_in_2968(dataIn[2968]),
.io_in_2969(dataIn[2969]),
.io_in_2970(dataIn[2970]),
.io_in_2971(dataIn[2971]),
.io_in_2972(dataIn[2972]),
.io_in_2973(dataIn[2973]),
.io_in_2974(dataIn[2974]),
.io_in_2975(dataIn[2975]),
.io_in_2976(dataIn[2976]),
.io_in_2977(dataIn[2977]),
.io_in_2978(dataIn[2978]),
.io_in_2979(dataIn[2979]),
.io_in_2980(dataIn[2980]),
.io_in_2981(dataIn[2981]),
.io_in_2982(dataIn[2982]),
.io_in_2983(dataIn[2983]),
.io_in_2984(dataIn[2984]),
.io_in_2985(dataIn[2985]),
.io_in_2986(dataIn[2986]),
.io_in_2987(dataIn[2987]),
.io_in_2988(dataIn[2988]),
.io_in_2989(dataIn[2989]),
.io_in_2990(dataIn[2990]),
.io_in_2991(dataIn[2991]),
.io_in_2992(dataIn[2992]),
.io_in_2993(dataIn[2993]),
.io_in_2994(dataIn[2994]),
.io_in_2995(dataIn[2995]),
.io_in_2996(dataIn[2996]),
.io_in_2997(dataIn[2997]),
.io_in_2998(dataIn[2998]),
.io_in_2999(dataIn[2999]),
.io_in_3000(dataIn[3000]),
.io_in_3001(dataIn[3001]),
.io_in_3002(dataIn[3002]),
.io_in_3003(dataIn[3003]),
.io_in_3004(dataIn[3004]),
.io_in_3005(dataIn[3005]),
.io_in_3006(dataIn[3006]),
.io_in_3007(dataIn[3007]),
.io_in_3008(dataIn[3008]),
.io_in_3009(dataIn[3009]),
.io_in_3010(dataIn[3010]),
.io_in_3011(dataIn[3011]),
.io_in_3012(dataIn[3012]),
.io_in_3013(dataIn[3013]),
.io_in_3014(dataIn[3014]),
.io_in_3015(dataIn[3015]),
.io_in_3016(dataIn[3016]),
.io_in_3017(dataIn[3017]),
.io_in_3018(dataIn[3018]),
.io_in_3019(dataIn[3019]),
.io_in_3020(dataIn[3020]),
.io_in_3021(dataIn[3021]),
.io_in_3022(dataIn[3022]),
.io_in_3023(dataIn[3023]),
.io_in_3024(dataIn[3024]),
.io_in_3025(dataIn[3025]),
.io_in_3026(dataIn[3026]),
.io_in_3027(dataIn[3027]),
.io_in_3028(dataIn[3028]),
.io_in_3029(dataIn[3029]),
.io_in_3030(dataIn[3030]),
.io_in_3031(dataIn[3031]),
.io_in_3032(dataIn[3032]),
.io_in_3033(dataIn[3033]),
.io_in_3034(dataIn[3034]),
.io_in_3035(dataIn[3035]),
.io_in_3036(dataIn[3036]),
.io_in_3037(dataIn[3037]),
.io_in_3038(dataIn[3038]),
.io_in_3039(dataIn[3039]),
.io_in_3040(dataIn[3040]),
.io_in_3041(dataIn[3041]),
.io_in_3042(dataIn[3042]),
.io_in_3043(dataIn[3043]),
.io_in_3044(dataIn[3044]),
.io_in_3045(dataIn[3045]),
.io_in_3046(dataIn[3046]),
.io_in_3047(dataIn[3047]),
.io_in_3048(dataIn[3048]),
.io_in_3049(dataIn[3049]),
.io_in_3050(dataIn[3050]),
.io_in_3051(dataIn[3051]),
.io_in_3052(dataIn[3052]),
.io_in_3053(dataIn[3053]),
.io_in_3054(dataIn[3054]),
.io_in_3055(dataIn[3055]),
.io_in_3056(dataIn[3056]),
.io_in_3057(dataIn[3057]),
.io_in_3058(dataIn[3058]),
.io_in_3059(dataIn[3059]),
.io_in_3060(dataIn[3060]),
.io_in_3061(dataIn[3061]),
.io_in_3062(dataIn[3062]),
.io_in_3063(dataIn[3063]),
.io_in_3064(dataIn[3064]),
.io_in_3065(dataIn[3065]),
.io_in_3066(dataIn[3066]),
.io_in_3067(dataIn[3067]),
.io_in_3068(dataIn[3068]),
.io_in_3069(dataIn[3069]),
.io_in_3070(dataIn[3070]),
.io_in_3071(dataIn[3071]),
.io_in_3072(dataIn[3072]),
.io_in_3073(dataIn[3073]),
.io_in_3074(dataIn[3074]),
.io_in_3075(dataIn[3075]),
.io_in_3076(dataIn[3076]),
.io_in_3077(dataIn[3077]),
.io_in_3078(dataIn[3078]),
.io_in_3079(dataIn[3079]),
.io_in_3080(dataIn[3080]),
.io_in_3081(dataIn[3081]),
.io_in_3082(dataIn[3082]),
.io_in_3083(dataIn[3083]),
.io_in_3084(dataIn[3084]),
.io_in_3085(dataIn[3085]),
.io_in_3086(dataIn[3086]),
.io_in_3087(dataIn[3087]),
.io_in_3088(dataIn[3088]),
.io_in_3089(dataIn[3089]),
.io_in_3090(dataIn[3090]),
.io_in_3091(dataIn[3091]),
.io_in_3092(dataIn[3092]),
.io_in_3093(dataIn[3093]),
.io_in_3094(dataIn[3094]),
.io_in_3095(dataIn[3095]),
.io_in_3096(dataIn[3096]),
.io_in_3097(dataIn[3097]),
.io_in_3098(dataIn[3098]),
.io_in_3099(dataIn[3099]),
.io_in_3100(dataIn[3100]),
.io_in_3101(dataIn[3101]),
.io_in_3102(dataIn[3102]),
.io_in_3103(dataIn[3103]),
.io_in_3104(dataIn[3104]),
.io_in_3105(dataIn[3105]),
.io_in_3106(dataIn[3106]),
.io_in_3107(dataIn[3107]),
.io_in_3108(dataIn[3108]),
.io_in_3109(dataIn[3109]),
.io_in_3110(dataIn[3110]),
.io_in_3111(dataIn[3111]),
.io_in_3112(dataIn[3112]),
.io_in_3113(dataIn[3113]),
.io_in_3114(dataIn[3114]),
.io_in_3115(dataIn[3115]),
.io_in_3116(dataIn[3116]),
.io_in_3117(dataIn[3117]),
.io_in_3118(dataIn[3118]),
.io_in_3119(dataIn[3119]),
.io_in_3120(dataIn[3120]),
.io_in_3121(dataIn[3121]),
.io_in_3122(dataIn[3122]),
.io_in_3123(dataIn[3123]),
.io_in_3124(dataIn[3124]),
.io_in_3125(dataIn[3125]),
.io_in_3126(dataIn[3126]),
.io_in_3127(dataIn[3127]),
.io_in_3128(dataIn[3128]),
.io_in_3129(dataIn[3129]),
.io_in_3130(dataIn[3130]),
.io_in_3131(dataIn[3131]),
.io_in_3132(dataIn[3132]),
.io_in_3133(dataIn[3133]),
.io_in_3134(dataIn[3134]),
.io_in_3135(dataIn[3135]),
.io_in_3136(dataIn[3136]),
.io_in_3137(dataIn[3137]),
.io_in_3138(dataIn[3138]),
.io_in_3139(dataIn[3139]),
.io_in_3140(dataIn[3140]),
.io_in_3141(dataIn[3141]),
.io_in_3142(dataIn[3142]),
.io_in_3143(dataIn[3143]),
.io_in_3144(dataIn[3144]),
.io_in_3145(dataIn[3145]),
.io_in_3146(dataIn[3146]),
.io_in_3147(dataIn[3147]),
.io_in_3148(dataIn[3148]),
.io_in_3149(dataIn[3149]),
.io_in_3150(dataIn[3150]),
.io_in_3151(dataIn[3151]),
.io_in_3152(dataIn[3152]),
.io_in_3153(dataIn[3153]),
.io_in_3154(dataIn[3154]),
.io_in_3155(dataIn[3155]),
.io_in_3156(dataIn[3156]),
.io_in_3157(dataIn[3157]),
.io_in_3158(dataIn[3158]),
.io_in_3159(dataIn[3159]),
.io_in_3160(dataIn[3160]),
.io_in_3161(dataIn[3161]),
.io_in_3162(dataIn[3162]),
.io_in_3163(dataIn[3163]),
.io_in_3164(dataIn[3164]),
.io_in_3165(dataIn[3165]),
.io_in_3166(dataIn[3166]),
.io_in_3167(dataIn[3167]),
.io_in_3168(dataIn[3168]),
.io_in_3169(dataIn[3169]),
.io_in_3170(dataIn[3170]),
.io_in_3171(dataIn[3171]),
.io_in_3172(dataIn[3172]),
.io_in_3173(dataIn[3173]),
.io_in_3174(dataIn[3174]),
.io_in_3175(dataIn[3175]),
.io_in_3176(dataIn[3176]),
.io_in_3177(dataIn[3177]),
.io_in_3178(dataIn[3178]),
.io_in_3179(dataIn[3179]),
.io_in_3180(dataIn[3180]),
.io_in_3181(dataIn[3181]),
.io_in_3182(dataIn[3182]),
.io_in_3183(dataIn[3183]),
.io_in_3184(dataIn[3184]),
.io_in_3185(dataIn[3185]),
.io_in_3186(dataIn[3186]),
.io_in_3187(dataIn[3187]),
.io_in_3188(dataIn[3188]),
.io_in_3189(dataIn[3189]),
.io_in_3190(dataIn[3190]),
.io_in_3191(dataIn[3191]),
.io_in_3192(dataIn[3192]),
.io_in_3193(dataIn[3193]),
.io_in_3194(dataIn[3194]),
.io_in_3195(dataIn[3195]),
.io_in_3196(dataIn[3196]),
.io_in_3197(dataIn[3197]),
.io_in_3198(dataIn[3198]),
.io_in_3199(dataIn[3199]),
.io_in_3200(dataIn[3200]),
.io_in_3201(dataIn[3201]),
.io_in_3202(dataIn[3202]),
.io_in_3203(dataIn[3203]),
.io_in_3204(dataIn[3204]),
.io_in_3205(dataIn[3205]),
.io_in_3206(dataIn[3206]),
.io_in_3207(dataIn[3207]),
.io_in_3208(dataIn[3208]),
.io_in_3209(dataIn[3209]),
.io_in_3210(dataIn[3210]),
.io_in_3211(dataIn[3211]),
.io_in_3212(dataIn[3212]),
.io_in_3213(dataIn[3213]),
.io_in_3214(dataIn[3214]),
.io_in_3215(dataIn[3215]),
.io_in_3216(dataIn[3216]),
.io_in_3217(dataIn[3217]),
.io_in_3218(dataIn[3218]),
.io_in_3219(dataIn[3219]),
.io_in_3220(dataIn[3220]),
.io_in_3221(dataIn[3221]),
.io_in_3222(dataIn[3222]),
.io_in_3223(dataIn[3223]),
.io_in_3224(dataIn[3224]),
.io_in_3225(dataIn[3225]),
.io_in_3226(dataIn[3226]),
.io_in_3227(dataIn[3227]),
.io_in_3228(dataIn[3228]),
.io_in_3229(dataIn[3229]),
.io_in_3230(dataIn[3230]),
.io_in_3231(dataIn[3231]),
.io_in_3232(dataIn[3232]),
.io_in_3233(dataIn[3233]),
.io_in_3234(dataIn[3234]),
.io_in_3235(dataIn[3235]),
.io_in_3236(dataIn[3236]),
.io_in_3237(dataIn[3237]),
.io_in_3238(dataIn[3238]),
.io_in_3239(dataIn[3239]),
.io_in_3240(dataIn[3240]),
.io_in_3241(dataIn[3241]),
.io_in_3242(dataIn[3242]),
.io_in_3243(dataIn[3243]),
.io_in_3244(dataIn[3244]),
.io_in_3245(dataIn[3245]),
.io_in_3246(dataIn[3246]),
.io_in_3247(dataIn[3247]),
.io_in_3248(dataIn[3248]),
.io_in_3249(dataIn[3249]),
.io_in_3250(dataIn[3250]),
.io_in_3251(dataIn[3251]),
.io_in_3252(dataIn[3252]),
.io_in_3253(dataIn[3253]),
.io_in_3254(dataIn[3254]),
.io_in_3255(dataIn[3255]),
.io_in_3256(dataIn[3256]),
.io_in_3257(dataIn[3257]),
.io_in_3258(dataIn[3258]),
.io_in_3259(dataIn[3259]),
.io_in_3260(dataIn[3260]),
.io_in_3261(dataIn[3261]),
.io_in_3262(dataIn[3262]),
.io_in_3263(dataIn[3263]),
.io_in_3264(dataIn[3264]),
.io_in_3265(dataIn[3265]),
.io_in_3266(dataIn[3266]),
.io_in_3267(dataIn[3267]),
.io_in_3268(dataIn[3268]),
.io_in_3269(dataIn[3269]),
.io_in_3270(dataIn[3270]),
.io_in_3271(dataIn[3271]),
.io_in_3272(dataIn[3272]),
.io_in_3273(dataIn[3273]),
.io_in_3274(dataIn[3274]),
.io_in_3275(dataIn[3275]),
.io_in_3276(dataIn[3276]),
.io_in_3277(dataIn[3277]),
.io_in_3278(dataIn[3278]),
.io_in_3279(dataIn[3279]),
.io_in_3280(dataIn[3280]),
.io_in_3281(dataIn[3281]),
.io_in_3282(dataIn[3282]),
.io_in_3283(dataIn[3283]),
.io_in_3284(dataIn[3284]),
.io_in_3285(dataIn[3285]),
.io_in_3286(dataIn[3286]),
.io_in_3287(dataIn[3287]),
.io_in_3288(dataIn[3288]),
.io_in_3289(dataIn[3289]),
.io_in_3290(dataIn[3290]),
.io_in_3291(dataIn[3291]),
.io_in_3292(dataIn[3292]),
.io_in_3293(dataIn[3293]),
.io_in_3294(dataIn[3294]),
.io_in_3295(dataIn[3295]),
.io_in_3296(dataIn[3296]),
.io_in_3297(dataIn[3297]),
.io_in_3298(dataIn[3298]),
.io_in_3299(dataIn[3299]),
.io_in_3300(dataIn[3300]),
.io_in_3301(dataIn[3301]),
.io_in_3302(dataIn[3302]),
.io_in_3303(dataIn[3303]),
.io_in_3304(dataIn[3304]),
.io_in_3305(dataIn[3305]),
.io_in_3306(dataIn[3306]),
.io_in_3307(dataIn[3307]),
.io_in_3308(dataIn[3308]),
.io_in_3309(dataIn[3309]),
.io_in_3310(dataIn[3310]),
.io_in_3311(dataIn[3311]),
.io_in_3312(dataIn[3312]),
.io_in_3313(dataIn[3313]),
.io_in_3314(dataIn[3314]),
.io_in_3315(dataIn[3315]),
.io_in_3316(dataIn[3316]),
.io_in_3317(dataIn[3317]),
.io_in_3318(dataIn[3318]),
.io_in_3319(dataIn[3319]),
.io_in_3320(dataIn[3320]),
.io_in_3321(dataIn[3321]),
.io_in_3322(dataIn[3322]),
.io_in_3323(dataIn[3323]),
.io_in_3324(dataIn[3324]),
.io_in_3325(dataIn[3325]),
.io_in_3326(dataIn[3326]),
.io_in_3327(dataIn[3327]),
.io_in_3328(dataIn[3328]),
.io_in_3329(dataIn[3329]),
.io_in_3330(dataIn[3330]),
.io_in_3331(dataIn[3331]),
.io_in_3332(dataIn[3332]),
.io_in_3333(dataIn[3333]),
.io_in_3334(dataIn[3334]),
.io_in_3335(dataIn[3335]),
.io_in_3336(dataIn[3336]),
.io_in_3337(dataIn[3337]),
.io_in_3338(dataIn[3338]),
.io_in_3339(dataIn[3339]),
.io_in_3340(dataIn[3340]),
.io_in_3341(dataIn[3341]),
.io_in_3342(dataIn[3342]),
.io_in_3343(dataIn[3343]),
.io_in_3344(dataIn[3344]),
.io_in_3345(dataIn[3345]),
.io_in_3346(dataIn[3346]),
.io_in_3347(dataIn[3347]),
.io_in_3348(dataIn[3348]),
.io_in_3349(dataIn[3349]),
.io_in_3350(dataIn[3350]),
.io_in_3351(dataIn[3351]),
.io_in_3352(dataIn[3352]),
.io_in_3353(dataIn[3353]),
.io_in_3354(dataIn[3354]),
.io_in_3355(dataIn[3355]),
.io_in_3356(dataIn[3356]),
.io_in_3357(dataIn[3357]),
.io_in_3358(dataIn[3358]),
.io_in_3359(dataIn[3359]),
.io_in_3360(dataIn[3360]),
.io_in_3361(dataIn[3361]),
.io_in_3362(dataIn[3362]),
.io_in_3363(dataIn[3363]),
.io_in_3364(dataIn[3364]),
.io_in_3365(dataIn[3365]),
.io_in_3366(dataIn[3366]),
.io_in_3367(dataIn[3367]),
.io_in_3368(dataIn[3368]),
.io_in_3369(dataIn[3369]),
.io_in_3370(dataIn[3370]),
.io_in_3371(dataIn[3371]),
.io_in_3372(dataIn[3372]),
.io_in_3373(dataIn[3373]),
.io_in_3374(dataIn[3374]),
.io_in_3375(dataIn[3375]),
.io_in_3376(dataIn[3376]),
.io_in_3377(dataIn[3377]),
.io_in_3378(dataIn[3378]),
.io_in_3379(dataIn[3379]),
.io_in_3380(dataIn[3380]),
.io_in_3381(dataIn[3381]),
.io_in_3382(dataIn[3382]),
.io_in_3383(dataIn[3383]),
.io_in_3384(dataIn[3384]),
.io_in_3385(dataIn[3385]),
.io_in_3386(dataIn[3386]),
.io_in_3387(dataIn[3387]),
.io_in_3388(dataIn[3388]),
.io_in_3389(dataIn[3389]),
.io_in_3390(dataIn[3390]),
.io_in_3391(dataIn[3391]),
.io_in_3392(dataIn[3392]),
.io_in_3393(dataIn[3393]),
.io_in_3394(dataIn[3394]),
.io_in_3395(dataIn[3395]),
.io_in_3396(dataIn[3396]),
.io_in_3397(dataIn[3397]),
.io_in_3398(dataIn[3398]),
.io_in_3399(dataIn[3399]),
.io_in_3400(dataIn[3400]),
.io_in_3401(dataIn[3401]),
.io_in_3402(dataIn[3402]),
.io_in_3403(dataIn[3403]),
.io_in_3404(dataIn[3404]),
.io_in_3405(dataIn[3405]),
.io_in_3406(dataIn[3406]),
.io_in_3407(dataIn[3407]),
.io_in_3408(dataIn[3408]),
.io_in_3409(dataIn[3409]),
.io_in_3410(dataIn[3410]),
.io_in_3411(dataIn[3411]),
.io_in_3412(dataIn[3412]),
.io_in_3413(dataIn[3413]),
.io_in_3414(dataIn[3414]),
.io_in_3415(dataIn[3415]),
.io_in_3416(dataIn[3416]),
.io_in_3417(dataIn[3417]),
.io_in_3418(dataIn[3418]),
.io_in_3419(dataIn[3419]),
.io_in_3420(dataIn[3420]),
.io_in_3421(dataIn[3421]),
.io_in_3422(dataIn[3422]),
.io_in_3423(dataIn[3423]),
.io_in_3424(dataIn[3424]),
.io_in_3425(dataIn[3425]),
.io_in_3426(dataIn[3426]),
.io_in_3427(dataIn[3427]),
.io_in_3428(dataIn[3428]),
.io_in_3429(dataIn[3429]),
.io_in_3430(dataIn[3430]),
.io_in_3431(dataIn[3431]),
.io_in_3432(dataIn[3432]),
.io_in_3433(dataIn[3433]),
.io_in_3434(dataIn[3434]),
.io_in_3435(dataIn[3435]),
.io_in_3436(dataIn[3436]),
.io_in_3437(dataIn[3437]),
.io_in_3438(dataIn[3438]),
.io_in_3439(dataIn[3439]),
.io_in_3440(dataIn[3440]),
.io_in_3441(dataIn[3441]),
.io_in_3442(dataIn[3442]),
.io_in_3443(dataIn[3443]),
.io_in_3444(dataIn[3444]),
.io_in_3445(dataIn[3445]),
.io_in_3446(dataIn[3446]),
.io_in_3447(dataIn[3447]),
.io_in_3448(dataIn[3448]),
.io_in_3449(dataIn[3449]),
.io_in_3450(dataIn[3450]),
.io_in_3451(dataIn[3451]),
.io_in_3452(dataIn[3452]),
.io_in_3453(dataIn[3453]),
.io_in_3454(dataIn[3454]),
.io_in_3455(dataIn[3455]),
.io_in_3456(dataIn[3456]),
.io_in_3457(dataIn[3457]),
.io_in_3458(dataIn[3458]),
.io_in_3459(dataIn[3459]),
.io_in_3460(dataIn[3460]),
.io_in_3461(dataIn[3461]),
.io_in_3462(dataIn[3462]),
.io_in_3463(dataIn[3463]),
.io_in_3464(dataIn[3464]),
.io_in_3465(dataIn[3465]),
.io_in_3466(dataIn[3466]),
.io_in_3467(dataIn[3467]),
.io_in_3468(dataIn[3468]),
.io_in_3469(dataIn[3469]),
.io_in_3470(dataIn[3470]),
.io_in_3471(dataIn[3471]),
.io_in_3472(dataIn[3472]),
.io_in_3473(dataIn[3473]),
.io_in_3474(dataIn[3474]),
.io_in_3475(dataIn[3475]),
.io_in_3476(dataIn[3476]),
.io_in_3477(dataIn[3477]),
.io_in_3478(dataIn[3478]),
.io_in_3479(dataIn[3479]),
.io_in_3480(dataIn[3480]),
.io_in_3481(dataIn[3481]),
.io_in_3482(dataIn[3482]),
.io_in_3483(dataIn[3483]),
.io_in_3484(dataIn[3484]),
.io_in_3485(dataIn[3485]),
.io_in_3486(dataIn[3486]),
.io_in_3487(dataIn[3487]),
.io_in_3488(dataIn[3488]),
.io_in_3489(dataIn[3489]),
.io_in_3490(dataIn[3490]),
.io_in_3491(dataIn[3491]),
.io_in_3492(dataIn[3492]),
.io_in_3493(dataIn[3493]),
.io_in_3494(dataIn[3494]),
.io_in_3495(dataIn[3495]),
.io_in_3496(dataIn[3496]),
.io_in_3497(dataIn[3497]),
.io_in_3498(dataIn[3498]),
.io_in_3499(dataIn[3499]),
.io_in_3500(dataIn[3500]),
.io_in_3501(dataIn[3501]),
.io_in_3502(dataIn[3502]),
.io_in_3503(dataIn[3503]),
.io_in_3504(dataIn[3504]),
.io_in_3505(dataIn[3505]),
.io_in_3506(dataIn[3506]),
.io_in_3507(dataIn[3507]),
.io_in_3508(dataIn[3508]),
.io_in_3509(dataIn[3509]),
.io_in_3510(dataIn[3510]),
.io_in_3511(dataIn[3511]),
.io_in_3512(dataIn[3512]),
.io_in_3513(dataIn[3513]),
.io_in_3514(dataIn[3514]),
.io_in_3515(dataIn[3515]),
.io_in_3516(dataIn[3516]),
.io_in_3517(dataIn[3517]),
.io_in_3518(dataIn[3518]),
.io_in_3519(dataIn[3519]),
.io_in_3520(dataIn[3520]),
.io_in_3521(dataIn[3521]),
.io_in_3522(dataIn[3522]),
.io_in_3523(dataIn[3523]),
.io_in_3524(dataIn[3524]),
.io_in_3525(dataIn[3525]),
.io_in_3526(dataIn[3526]),
.io_in_3527(dataIn[3527]),
.io_in_3528(dataIn[3528]),
.io_in_3529(dataIn[3529]),
.io_in_3530(dataIn[3530]),
.io_in_3531(dataIn[3531]),
.io_in_3532(dataIn[3532]),
.io_in_3533(dataIn[3533]),
.io_in_3534(dataIn[3534]),
.io_in_3535(dataIn[3535]),
.io_in_3536(dataIn[3536]),
.io_in_3537(dataIn[3537]),
.io_in_3538(dataIn[3538]),
.io_in_3539(dataIn[3539]),
.io_in_3540(dataIn[3540]),
.io_in_3541(dataIn[3541]),
.io_in_3542(dataIn[3542]),
.io_in_3543(dataIn[3543]),
.io_in_3544(dataIn[3544]),
.io_in_3545(dataIn[3545]),
.io_in_3546(dataIn[3546]),
.io_in_3547(dataIn[3547]),
.io_in_3548(dataIn[3548]),
.io_in_3549(dataIn[3549]),
.io_in_3550(dataIn[3550]),
.io_in_3551(dataIn[3551]),
.io_in_3552(dataIn[3552]),
.io_in_3553(dataIn[3553]),
.io_in_3554(dataIn[3554]),
.io_in_3555(dataIn[3555]),
.io_in_3556(dataIn[3556]),
.io_in_3557(dataIn[3557]),
.io_in_3558(dataIn[3558]),
.io_in_3559(dataIn[3559]),
.io_in_3560(dataIn[3560]),
.io_in_3561(dataIn[3561]),
.io_in_3562(dataIn[3562]),
.io_in_3563(dataIn[3563]),
.io_in_3564(dataIn[3564]),
.io_in_3565(dataIn[3565]),
.io_in_3566(dataIn[3566]),
.io_in_3567(dataIn[3567]),
.io_in_3568(dataIn[3568]),
.io_in_3569(dataIn[3569]),
.io_in_3570(dataIn[3570]),
.io_in_3571(dataIn[3571]),
.io_in_3572(dataIn[3572]),
.io_in_3573(dataIn[3573]),
.io_in_3574(dataIn[3574]),
.io_in_3575(dataIn[3575]),
.io_in_3576(dataIn[3576]),
.io_in_3577(dataIn[3577]),
.io_in_3578(dataIn[3578]),
.io_in_3579(dataIn[3579]),
.io_in_3580(dataIn[3580]),
.io_in_3581(dataIn[3581]),
.io_in_3582(dataIn[3582]),
.io_in_3583(dataIn[3583]),
.io_in_3584(dataIn[3584]),
.io_in_3585(dataIn[3585]),
.io_in_3586(dataIn[3586]),
.io_in_3587(dataIn[3587]),
.io_in_3588(dataIn[3588]),
.io_in_3589(dataIn[3589]),
.io_in_3590(dataIn[3590]),
.io_in_3591(dataIn[3591]),
.io_in_3592(dataIn[3592]),
.io_in_3593(dataIn[3593]),
.io_in_3594(dataIn[3594]),
.io_in_3595(dataIn[3595]),
.io_in_3596(dataIn[3596]),
.io_in_3597(dataIn[3597]),
.io_in_3598(dataIn[3598]),
.io_in_3599(dataIn[3599]),
.io_in_3600(dataIn[3600]),
.io_in_3601(dataIn[3601]),
.io_in_3602(dataIn[3602]),
.io_in_3603(dataIn[3603]),
.io_in_3604(dataIn[3604]),
.io_in_3605(dataIn[3605]),
.io_in_3606(dataIn[3606]),
.io_in_3607(dataIn[3607]),
.io_in_3608(dataIn[3608]),
.io_in_3609(dataIn[3609]),
.io_in_3610(dataIn[3610]),
.io_in_3611(dataIn[3611]),
.io_in_3612(dataIn[3612]),
.io_in_3613(dataIn[3613]),
.io_in_3614(dataIn[3614]),
.io_in_3615(dataIn[3615]),
.io_in_3616(dataIn[3616]),
.io_in_3617(dataIn[3617]),
.io_in_3618(dataIn[3618]),
.io_in_3619(dataIn[3619]),
.io_in_3620(dataIn[3620]),
.io_in_3621(dataIn[3621]),
.io_in_3622(dataIn[3622]),
.io_in_3623(dataIn[3623]),
.io_in_3624(dataIn[3624]),
.io_in_3625(dataIn[3625]),
.io_in_3626(dataIn[3626]),
.io_in_3627(dataIn[3627]),
.io_in_3628(dataIn[3628]),
.io_in_3629(dataIn[3629]),
.io_in_3630(dataIn[3630]),
.io_in_3631(dataIn[3631]),
.io_in_3632(dataIn[3632]),
.io_in_3633(dataIn[3633]),
.io_in_3634(dataIn[3634]),
.io_in_3635(dataIn[3635]),
.io_in_3636(dataIn[3636]),
.io_in_3637(dataIn[3637]),
.io_in_3638(dataIn[3638]),
.io_in_3639(dataIn[3639]),
.io_in_3640(dataIn[3640]),
.io_in_3641(dataIn[3641]),
.io_in_3642(dataIn[3642]),
.io_in_3643(dataIn[3643]),
.io_in_3644(dataIn[3644]),
.io_in_3645(dataIn[3645]),
.io_in_3646(dataIn[3646]),
.io_in_3647(dataIn[3647]),
.io_in_3648(dataIn[3648]),
.io_in_3649(dataIn[3649]),
.io_in_3650(dataIn[3650]),
.io_in_3651(dataIn[3651]),
.io_in_3652(dataIn[3652]),
.io_in_3653(dataIn[3653]),
.io_in_3654(dataIn[3654]),
.io_in_3655(dataIn[3655]),
.io_in_3656(dataIn[3656]),
.io_in_3657(dataIn[3657]),
.io_in_3658(dataIn[3658]),
.io_in_3659(dataIn[3659]),
.io_in_3660(dataIn[3660]),
.io_in_3661(dataIn[3661]),
.io_in_3662(dataIn[3662]),
.io_in_3663(dataIn[3663]),
.io_in_3664(dataIn[3664]),
.io_in_3665(dataIn[3665]),
.io_in_3666(dataIn[3666]),
.io_in_3667(dataIn[3667]),
.io_in_3668(dataIn[3668]),
.io_in_3669(dataIn[3669]),
.io_in_3670(dataIn[3670]),
.io_in_3671(dataIn[3671]),
.io_in_3672(dataIn[3672]),
.io_in_3673(dataIn[3673]),
.io_in_3674(dataIn[3674]),
.io_in_3675(dataIn[3675]),
.io_in_3676(dataIn[3676]),
.io_in_3677(dataIn[3677]),
.io_in_3678(dataIn[3678]),
.io_in_3679(dataIn[3679]),
.io_in_3680(dataIn[3680]),
.io_in_3681(dataIn[3681]),
.io_in_3682(dataIn[3682]),
.io_in_3683(dataIn[3683]),
.io_in_3684(dataIn[3684]),
.io_in_3685(dataIn[3685]),
.io_in_3686(dataIn[3686]),
.io_in_3687(dataIn[3687]),
.io_in_3688(dataIn[3688]),
.io_in_3689(dataIn[3689]),
.io_in_3690(dataIn[3690]),
.io_in_3691(dataIn[3691]),
.io_in_3692(dataIn[3692]),
.io_in_3693(dataIn[3693]),
.io_in_3694(dataIn[3694]),
.io_in_3695(dataIn[3695]),
.io_in_3696(dataIn[3696]),
.io_in_3697(dataIn[3697]),
.io_in_3698(dataIn[3698]),
.io_in_3699(dataIn[3699]),
.io_in_3700(dataIn[3700]),
.io_in_3701(dataIn[3701]),
.io_in_3702(dataIn[3702]),
.io_in_3703(dataIn[3703]),
.io_in_3704(dataIn[3704]),
.io_in_3705(dataIn[3705]),
.io_in_3706(dataIn[3706]),
.io_in_3707(dataIn[3707]),
.io_in_3708(dataIn[3708]),
.io_in_3709(dataIn[3709]),
.io_in_3710(dataIn[3710]),
.io_in_3711(dataIn[3711]),
.io_in_3712(dataIn[3712]),
.io_in_3713(dataIn[3713]),
.io_in_3714(dataIn[3714]),
.io_in_3715(dataIn[3715]),
.io_in_3716(dataIn[3716]),
.io_in_3717(dataIn[3717]),
.io_in_3718(dataIn[3718]),
.io_in_3719(dataIn[3719]),
.io_in_3720(dataIn[3720]),
.io_in_3721(dataIn[3721]),
.io_in_3722(dataIn[3722]),
.io_in_3723(dataIn[3723]),
.io_in_3724(dataIn[3724]),
.io_in_3725(dataIn[3725]),
.io_in_3726(dataIn[3726]),
.io_in_3727(dataIn[3727]),
.io_in_3728(dataIn[3728]),
.io_in_3729(dataIn[3729]),
.io_in_3730(dataIn[3730]),
.io_in_3731(dataIn[3731]),
.io_in_3732(dataIn[3732]),
.io_in_3733(dataIn[3733]),
.io_in_3734(dataIn[3734]),
.io_in_3735(dataIn[3735]),
.io_in_3736(dataIn[3736]),
.io_in_3737(dataIn[3737]),
.io_in_3738(dataIn[3738]),
.io_in_3739(dataIn[3739]),
.io_in_3740(dataIn[3740]),
.io_in_3741(dataIn[3741]),
.io_in_3742(dataIn[3742]),
.io_in_3743(dataIn[3743]),
.io_in_3744(dataIn[3744]),
.io_in_3745(dataIn[3745]),
.io_in_3746(dataIn[3746]),
.io_in_3747(dataIn[3747]),
.io_in_3748(dataIn[3748]),
.io_in_3749(dataIn[3749]),
.io_in_3750(dataIn[3750]),
.io_in_3751(dataIn[3751]),
.io_in_3752(dataIn[3752]),
.io_in_3753(dataIn[3753]),
.io_in_3754(dataIn[3754]),
.io_in_3755(dataIn[3755]),
.io_in_3756(dataIn[3756]),
.io_in_3757(dataIn[3757]),
.io_in_3758(dataIn[3758]),
.io_in_3759(dataIn[3759]),
.io_in_3760(dataIn[3760]),
.io_in_3761(dataIn[3761]),
.io_in_3762(dataIn[3762]),
.io_in_3763(dataIn[3763]),
.io_in_3764(dataIn[3764]),
.io_in_3765(dataIn[3765]),
.io_in_3766(dataIn[3766]),
.io_in_3767(dataIn[3767]),
.io_in_3768(dataIn[3768]),
.io_in_3769(dataIn[3769]),
.io_in_3770(dataIn[3770]),
.io_in_3771(dataIn[3771]),
.io_in_3772(dataIn[3772]),
.io_in_3773(dataIn[3773]),
.io_in_3774(dataIn[3774]),
.io_in_3775(dataIn[3775]),
.io_in_3776(dataIn[3776]),
.io_in_3777(dataIn[3777]),
.io_in_3778(dataIn[3778]),
.io_in_3779(dataIn[3779]),
.io_in_3780(dataIn[3780]),
.io_in_3781(dataIn[3781]),
.io_in_3782(dataIn[3782]),
.io_in_3783(dataIn[3783]),
.io_in_3784(dataIn[3784]),
.io_in_3785(dataIn[3785]),
.io_in_3786(dataIn[3786]),
.io_in_3787(dataIn[3787]),
.io_in_3788(dataIn[3788]),
.io_in_3789(dataIn[3789]),
.io_in_3790(dataIn[3790]),
.io_in_3791(dataIn[3791]),
.io_in_3792(dataIn[3792]),
.io_in_3793(dataIn[3793]),
.io_in_3794(dataIn[3794]),
.io_in_3795(dataIn[3795]),
.io_in_3796(dataIn[3796]),
.io_in_3797(dataIn[3797]),
.io_in_3798(dataIn[3798]),
.io_in_3799(dataIn[3799]),
.io_in_3800(dataIn[3800]),
.io_in_3801(dataIn[3801]),
.io_in_3802(dataIn[3802]),
.io_in_3803(dataIn[3803]),
.io_in_3804(dataIn[3804]),
.io_in_3805(dataIn[3805]),
.io_in_3806(dataIn[3806]),
.io_in_3807(dataIn[3807]),
.io_in_3808(dataIn[3808]),
.io_in_3809(dataIn[3809]),
.io_in_3810(dataIn[3810]),
.io_in_3811(dataIn[3811]),
.io_in_3812(dataIn[3812]),
.io_in_3813(dataIn[3813]),
.io_in_3814(dataIn[3814]),
.io_in_3815(dataIn[3815]),
.io_in_3816(dataIn[3816]),
.io_in_3817(dataIn[3817]),
.io_in_3818(dataIn[3818]),
.io_in_3819(dataIn[3819]),
.io_in_3820(dataIn[3820]),
.io_in_3821(dataIn[3821]),
.io_in_3822(dataIn[3822]),
.io_in_3823(dataIn[3823]),
.io_in_3824(dataIn[3824]),
.io_in_3825(dataIn[3825]),
.io_in_3826(dataIn[3826]),
.io_in_3827(dataIn[3827]),
.io_in_3828(dataIn[3828]),
.io_in_3829(dataIn[3829]),
.io_in_3830(dataIn[3830]),
.io_in_3831(dataIn[3831]),
.io_in_3832(dataIn[3832]),
.io_in_3833(dataIn[3833]),
.io_in_3834(dataIn[3834]),
.io_in_3835(dataIn[3835]),
.io_in_3836(dataIn[3836]),
.io_in_3837(dataIn[3837]),
.io_in_3838(dataIn[3838]),
.io_in_3839(dataIn[3839]),
.io_in_3840(dataIn[3840]),
.io_in_3841(dataIn[3841]),
.io_in_3842(dataIn[3842]),
.io_in_3843(dataIn[3843]),
.io_in_3844(dataIn[3844]),
.io_in_3845(dataIn[3845]),
.io_in_3846(dataIn[3846]),
.io_in_3847(dataIn[3847]),
.io_in_3848(dataIn[3848]),
.io_in_3849(dataIn[3849]),
.io_in_3850(dataIn[3850]),
.io_in_3851(dataIn[3851]),
.io_in_3852(dataIn[3852]),
.io_in_3853(dataIn[3853]),
.io_in_3854(dataIn[3854]),
.io_in_3855(dataIn[3855]),
.io_in_3856(dataIn[3856]),
.io_in_3857(dataIn[3857]),
.io_in_3858(dataIn[3858]),
.io_in_3859(dataIn[3859]),
.io_in_3860(dataIn[3860]),
.io_in_3861(dataIn[3861]),
.io_in_3862(dataIn[3862]),
.io_in_3863(dataIn[3863]),
.io_in_3864(dataIn[3864]),
.io_in_3865(dataIn[3865]),
.io_in_3866(dataIn[3866]),
.io_in_3867(dataIn[3867]),
.io_in_3868(dataIn[3868]),
.io_in_3869(dataIn[3869]),
.io_in_3870(dataIn[3870]),
.io_in_3871(dataIn[3871]),
.io_in_3872(dataIn[3872]),
.io_in_3873(dataIn[3873]),
.io_in_3874(dataIn[3874]),
.io_in_3875(dataIn[3875]),
.io_in_3876(dataIn[3876]),
.io_in_3877(dataIn[3877]),
.io_in_3878(dataIn[3878]),
.io_in_3879(dataIn[3879]),
.io_in_3880(dataIn[3880]),
.io_in_3881(dataIn[3881]),
.io_in_3882(dataIn[3882]),
.io_in_3883(dataIn[3883]),
.io_in_3884(dataIn[3884]),
.io_in_3885(dataIn[3885]),
.io_in_3886(dataIn[3886]),
.io_in_3887(dataIn[3887]),
.io_in_3888(dataIn[3888]),
.io_in_3889(dataIn[3889]),
.io_in_3890(dataIn[3890]),
.io_in_3891(dataIn[3891]),
.io_in_3892(dataIn[3892]),
.io_in_3893(dataIn[3893]),
.io_in_3894(dataIn[3894]),
.io_in_3895(dataIn[3895]),
.io_in_3896(dataIn[3896]),
.io_in_3897(dataIn[3897]),
.io_in_3898(dataIn[3898]),
.io_in_3899(dataIn[3899]),
.io_in_3900(dataIn[3900]),
.io_in_3901(dataIn[3901]),
.io_in_3902(dataIn[3902]),
.io_in_3903(dataIn[3903]),
.io_in_3904(dataIn[3904]),
.io_in_3905(dataIn[3905]),
.io_in_3906(dataIn[3906]),
.io_in_3907(dataIn[3907]),
.io_in_3908(dataIn[3908]),
.io_in_3909(dataIn[3909]),
.io_in_3910(dataIn[3910]),
.io_in_3911(dataIn[3911]),
.io_in_3912(dataIn[3912]),
.io_in_3913(dataIn[3913]),
.io_in_3914(dataIn[3914]),
.io_in_3915(dataIn[3915]),
.io_in_3916(dataIn[3916]),
.io_in_3917(dataIn[3917]),
.io_in_3918(dataIn[3918]),
.io_in_3919(dataIn[3919]),
.io_in_3920(dataIn[3920]),
.io_in_3921(dataIn[3921]),
.io_in_3922(dataIn[3922]),
.io_in_3923(dataIn[3923]),
.io_in_3924(dataIn[3924]),
.io_in_3925(dataIn[3925]),
.io_in_3926(dataIn[3926]),
.io_in_3927(dataIn[3927]),
.io_in_3928(dataIn[3928]),
.io_in_3929(dataIn[3929]),
.io_in_3930(dataIn[3930]),
.io_in_3931(dataIn[3931]),
.io_in_3932(dataIn[3932]),
.io_in_3933(dataIn[3933]),
.io_in_3934(dataIn[3934]),
.io_in_3935(dataIn[3935]),
.io_in_3936(dataIn[3936]),
.io_in_3937(dataIn[3937]),
.io_in_3938(dataIn[3938]),
.io_in_3939(dataIn[3939]),
.io_in_3940(dataIn[3940]),
.io_in_3941(dataIn[3941]),
.io_in_3942(dataIn[3942]),
.io_in_3943(dataIn[3943]),
.io_in_3944(dataIn[3944]),
.io_in_3945(dataIn[3945]),
.io_in_3946(dataIn[3946]),
.io_in_3947(dataIn[3947]),
.io_in_3948(dataIn[3948]),
.io_in_3949(dataIn[3949]),
.io_in_3950(dataIn[3950]),
.io_in_3951(dataIn[3951]),
.io_in_3952(dataIn[3952]),
.io_in_3953(dataIn[3953]),
.io_in_3954(dataIn[3954]),
.io_in_3955(dataIn[3955]),
.io_in_3956(dataIn[3956]),
.io_in_3957(dataIn[3957]),
.io_in_3958(dataIn[3958]),
.io_in_3959(dataIn[3959]),
.io_in_3960(dataIn[3960]),
.io_in_3961(dataIn[3961]),
.io_in_3962(dataIn[3962]),
.io_in_3963(dataIn[3963]),
.io_in_3964(dataIn[3964]),
.io_in_3965(dataIn[3965]),
.io_in_3966(dataIn[3966]),
.io_in_3967(dataIn[3967]),
.io_in_3968(dataIn[3968]),
.io_in_3969(dataIn[3969]),
.io_in_3970(dataIn[3970]),
.io_in_3971(dataIn[3971]),
.io_in_3972(dataIn[3972]),
.io_in_3973(dataIn[3973]),
.io_in_3974(dataIn[3974]),
.io_in_3975(dataIn[3975]),
.io_in_3976(dataIn[3976]),
.io_in_3977(dataIn[3977]),
.io_in_3978(dataIn[3978]),
.io_in_3979(dataIn[3979]),
.io_in_3980(dataIn[3980]),
.io_in_3981(dataIn[3981]),
.io_in_3982(dataIn[3982]),
.io_in_3983(dataIn[3983]),
.io_in_3984(dataIn[3984]),
.io_in_3985(dataIn[3985]),
.io_in_3986(dataIn[3986]),
.io_in_3987(dataIn[3987]),
.io_in_3988(dataIn[3988]),
.io_in_3989(dataIn[3989]),
.io_in_3990(dataIn[3990]),
.io_in_3991(dataIn[3991]),
.io_in_3992(dataIn[3992]),
.io_in_3993(dataIn[3993]),
.io_in_3994(dataIn[3994]),
.io_in_3995(dataIn[3995]),
.io_in_3996(dataIn[3996]),
.io_in_3997(dataIn[3997]),
.io_in_3998(dataIn[3998]),
.io_in_3999(dataIn[3999]),
.io_in_4000(dataIn[4000]),
.io_in_4001(dataIn[4001]),
.io_in_4002(dataIn[4002]),
.io_in_4003(dataIn[4003]),
.io_in_4004(dataIn[4004]),
.io_in_4005(dataIn[4005]),
.io_in_4006(dataIn[4006]),
.io_in_4007(dataIn[4007]),
.io_in_4008(dataIn[4008]),
.io_in_4009(dataIn[4009]),
.io_in_4010(dataIn[4010]),
.io_in_4011(dataIn[4011]),
.io_in_4012(dataIn[4012]),
.io_in_4013(dataIn[4013]),
.io_in_4014(dataIn[4014]),
.io_in_4015(dataIn[4015]),
.io_in_4016(dataIn[4016]),
.io_in_4017(dataIn[4017]),
.io_in_4018(dataIn[4018]),
.io_in_4019(dataIn[4019]),
.io_in_4020(dataIn[4020]),
.io_in_4021(dataIn[4021]),
.io_in_4022(dataIn[4022]),
.io_in_4023(dataIn[4023]),
.io_in_4024(dataIn[4024]),
.io_in_4025(dataIn[4025]),
.io_in_4026(dataIn[4026]),
.io_in_4027(dataIn[4027]),
.io_in_4028(dataIn[4028]),
.io_in_4029(dataIn[4029]),
.io_in_4030(dataIn[4030]),
.io_in_4031(dataIn[4031]),
.io_in_4032(dataIn[4032]),
.io_in_4033(dataIn[4033]),
.io_in_4034(dataIn[4034]),
.io_in_4035(dataIn[4035]),
.io_in_4036(dataIn[4036]),
.io_in_4037(dataIn[4037]),
.io_in_4038(dataIn[4038]),
.io_in_4039(dataIn[4039]),
.io_in_4040(dataIn[4040]),
.io_in_4041(dataIn[4041]),
.io_in_4042(dataIn[4042]),
.io_in_4043(dataIn[4043]),
.io_in_4044(dataIn[4044]),
.io_in_4045(dataIn[4045]),
.io_in_4046(dataIn[4046]),
.io_in_4047(dataIn[4047]),
.io_in_4048(dataIn[4048]),
.io_in_4049(dataIn[4049]),
.io_in_4050(dataIn[4050]),
.io_in_4051(dataIn[4051]),
.io_in_4052(dataIn[4052]),
.io_in_4053(dataIn[4053]),
.io_in_4054(dataIn[4054]),
.io_in_4055(dataIn[4055]),
.io_in_4056(dataIn[4056]),
.io_in_4057(dataIn[4057]),
.io_in_4058(dataIn[4058]),
.io_in_4059(dataIn[4059]),
.io_in_4060(dataIn[4060]),
.io_in_4061(dataIn[4061]),
.io_in_4062(dataIn[4062]),
.io_in_4063(dataIn[4063]),
.io_in_4064(dataIn[4064]),
.io_in_4065(dataIn[4065]),
.io_in_4066(dataIn[4066]),
.io_in_4067(dataIn[4067]),
.io_in_4068(dataIn[4068]),
.io_in_4069(dataIn[4069]),
.io_in_4070(dataIn[4070]),
.io_in_4071(dataIn[4071]),
.io_in_4072(dataIn[4072]),
.io_in_4073(dataIn[4073]),
.io_in_4074(dataIn[4074]),
.io_in_4075(dataIn[4075]),
.io_in_4076(dataIn[4076]),
.io_in_4077(dataIn[4077]),
.io_in_4078(dataIn[4078]),
.io_in_4079(dataIn[4079]),
.io_in_4080(dataIn[4080]),
.io_in_4081(dataIn[4081]),
.io_in_4082(dataIn[4082]),
.io_in_4083(dataIn[4083]),
.io_in_4084(dataIn[4084]),
.io_in_4085(dataIn[4085]),
.io_in_4086(dataIn[4086]),
.io_in_4087(dataIn[4087]),
.io_in_4088(dataIn[4088]),
.io_in_4089(dataIn[4089]),
.io_in_4090(dataIn[4090]),
.io_in_4091(dataIn[4091]),
.io_in_4092(dataIn[4092]),
.io_in_4093(dataIn[4093]),
.io_in_4094(dataIn[4094]),
.io_in_4095(dataIn[4095]),
.io_out_0(dataOut[0]),
.io_out_1(dataOut[1]),
.io_out_2(dataOut[2]),
.io_out_3(dataOut[3]),
.io_out_4(dataOut[4]),
.io_out_5(dataOut[5]),
.io_out_6(dataOut[6]),
.io_out_7(dataOut[7]),
.io_out_8(dataOut[8]),
.io_out_9(dataOut[9]),
.io_out_10(dataOut[10]),
.io_out_11(dataOut[11]),
.io_out_12(dataOut[12]),
.io_out_13(dataOut[13]),
.io_out_14(dataOut[14]),
.io_out_15(dataOut[15]),
.io_out_16(dataOut[16]),
.io_out_17(dataOut[17]),
.io_out_18(dataOut[18]),
.io_out_19(dataOut[19]),
.io_out_20(dataOut[20]),
.io_out_21(dataOut[21]),
.io_out_22(dataOut[22]),
.io_out_23(dataOut[23]),
.io_out_24(dataOut[24]),
.io_out_25(dataOut[25]),
.io_out_26(dataOut[26]),
.io_out_27(dataOut[27]),
.io_out_28(dataOut[28]),
.io_out_29(dataOut[29]),
.io_out_30(dataOut[30]),
.io_out_31(dataOut[31]),
.io_out_32(dataOut[32]),
.io_out_33(dataOut[33]),
.io_out_34(dataOut[34]),
.io_out_35(dataOut[35]),
.io_out_36(dataOut[36]),
.io_out_37(dataOut[37]),
.io_out_38(dataOut[38]),
.io_out_39(dataOut[39]),
.io_out_40(dataOut[40]),
.io_out_41(dataOut[41]),
.io_out_42(dataOut[42]),
.io_out_43(dataOut[43]),
.io_out_44(dataOut[44]),
.io_out_45(dataOut[45]),
.io_out_46(dataOut[46]),
.io_out_47(dataOut[47]),
.io_out_48(dataOut[48]),
.io_out_49(dataOut[49]),
.io_out_50(dataOut[50]),
.io_out_51(dataOut[51]),
.io_out_52(dataOut[52]),
.io_out_53(dataOut[53]),
.io_out_54(dataOut[54]),
.io_out_55(dataOut[55]),
.io_out_56(dataOut[56]),
.io_out_57(dataOut[57]),
.io_out_58(dataOut[58]),
.io_out_59(dataOut[59]),
.io_out_60(dataOut[60]),
.io_out_61(dataOut[61]),
.io_out_62(dataOut[62]),
.io_out_63(dataOut[63]),
.io_out_64(dataOut[64]),
.io_out_65(dataOut[65]),
.io_out_66(dataOut[66]),
.io_out_67(dataOut[67]),
.io_out_68(dataOut[68]),
.io_out_69(dataOut[69]),
.io_out_70(dataOut[70]),
.io_out_71(dataOut[71]),
.io_out_72(dataOut[72]),
.io_out_73(dataOut[73]),
.io_out_74(dataOut[74]),
.io_out_75(dataOut[75]),
.io_out_76(dataOut[76]),
.io_out_77(dataOut[77]),
.io_out_78(dataOut[78]),
.io_out_79(dataOut[79]),
.io_out_80(dataOut[80]),
.io_out_81(dataOut[81]),
.io_out_82(dataOut[82]),
.io_out_83(dataOut[83]),
.io_out_84(dataOut[84]),
.io_out_85(dataOut[85]),
.io_out_86(dataOut[86]),
.io_out_87(dataOut[87]),
.io_out_88(dataOut[88]),
.io_out_89(dataOut[89]),
.io_out_90(dataOut[90]),
.io_out_91(dataOut[91]),
.io_out_92(dataOut[92]),
.io_out_93(dataOut[93]),
.io_out_94(dataOut[94]),
.io_out_95(dataOut[95]),
.io_out_96(dataOut[96]),
.io_out_97(dataOut[97]),
.io_out_98(dataOut[98]),
.io_out_99(dataOut[99]),
.io_out_100(dataOut[100]),
.io_out_101(dataOut[101]),
.io_out_102(dataOut[102]),
.io_out_103(dataOut[103]),
.io_out_104(dataOut[104]),
.io_out_105(dataOut[105]),
.io_out_106(dataOut[106]),
.io_out_107(dataOut[107]),
.io_out_108(dataOut[108]),
.io_out_109(dataOut[109]),
.io_out_110(dataOut[110]),
.io_out_111(dataOut[111]),
.io_out_112(dataOut[112]),
.io_out_113(dataOut[113]),
.io_out_114(dataOut[114]),
.io_out_115(dataOut[115]),
.io_out_116(dataOut[116]),
.io_out_117(dataOut[117]),
.io_out_118(dataOut[118]),
.io_out_119(dataOut[119]),
.io_out_120(dataOut[120]),
.io_out_121(dataOut[121]),
.io_out_122(dataOut[122]),
.io_out_123(dataOut[123]),
.io_out_124(dataOut[124]),
.io_out_125(dataOut[125]),
.io_out_126(dataOut[126]),
.io_out_127(dataOut[127]),
.io_out_128(dataOut[128]),
.io_out_129(dataOut[129]),
.io_out_130(dataOut[130]),
.io_out_131(dataOut[131]),
.io_out_132(dataOut[132]),
.io_out_133(dataOut[133]),
.io_out_134(dataOut[134]),
.io_out_135(dataOut[135]),
.io_out_136(dataOut[136]),
.io_out_137(dataOut[137]),
.io_out_138(dataOut[138]),
.io_out_139(dataOut[139]),
.io_out_140(dataOut[140]),
.io_out_141(dataOut[141]),
.io_out_142(dataOut[142]),
.io_out_143(dataOut[143]),
.io_out_144(dataOut[144]),
.io_out_145(dataOut[145]),
.io_out_146(dataOut[146]),
.io_out_147(dataOut[147]),
.io_out_148(dataOut[148]),
.io_out_149(dataOut[149]),
.io_out_150(dataOut[150]),
.io_out_151(dataOut[151]),
.io_out_152(dataOut[152]),
.io_out_153(dataOut[153]),
.io_out_154(dataOut[154]),
.io_out_155(dataOut[155]),
.io_out_156(dataOut[156]),
.io_out_157(dataOut[157]),
.io_out_158(dataOut[158]),
.io_out_159(dataOut[159]),
.io_out_160(dataOut[160]),
.io_out_161(dataOut[161]),
.io_out_162(dataOut[162]),
.io_out_163(dataOut[163]),
.io_out_164(dataOut[164]),
.io_out_165(dataOut[165]),
.io_out_166(dataOut[166]),
.io_out_167(dataOut[167]),
.io_out_168(dataOut[168]),
.io_out_169(dataOut[169]),
.io_out_170(dataOut[170]),
.io_out_171(dataOut[171]),
.io_out_172(dataOut[172]),
.io_out_173(dataOut[173]),
.io_out_174(dataOut[174]),
.io_out_175(dataOut[175]),
.io_out_176(dataOut[176]),
.io_out_177(dataOut[177]),
.io_out_178(dataOut[178]),
.io_out_179(dataOut[179]),
.io_out_180(dataOut[180]),
.io_out_181(dataOut[181]),
.io_out_182(dataOut[182]),
.io_out_183(dataOut[183]),
.io_out_184(dataOut[184]),
.io_out_185(dataOut[185]),
.io_out_186(dataOut[186]),
.io_out_187(dataOut[187]),
.io_out_188(dataOut[188]),
.io_out_189(dataOut[189]),
.io_out_190(dataOut[190]),
.io_out_191(dataOut[191]),
.io_out_192(dataOut[192]),
.io_out_193(dataOut[193]),
.io_out_194(dataOut[194]),
.io_out_195(dataOut[195]),
.io_out_196(dataOut[196]),
.io_out_197(dataOut[197]),
.io_out_198(dataOut[198]),
.io_out_199(dataOut[199]),
.io_out_200(dataOut[200]),
.io_out_201(dataOut[201]),
.io_out_202(dataOut[202]),
.io_out_203(dataOut[203]),
.io_out_204(dataOut[204]),
.io_out_205(dataOut[205]),
.io_out_206(dataOut[206]),
.io_out_207(dataOut[207]),
.io_out_208(dataOut[208]),
.io_out_209(dataOut[209]),
.io_out_210(dataOut[210]),
.io_out_211(dataOut[211]),
.io_out_212(dataOut[212]),
.io_out_213(dataOut[213]),
.io_out_214(dataOut[214]),
.io_out_215(dataOut[215]),
.io_out_216(dataOut[216]),
.io_out_217(dataOut[217]),
.io_out_218(dataOut[218]),
.io_out_219(dataOut[219]),
.io_out_220(dataOut[220]),
.io_out_221(dataOut[221]),
.io_out_222(dataOut[222]),
.io_out_223(dataOut[223]),
.io_out_224(dataOut[224]),
.io_out_225(dataOut[225]),
.io_out_226(dataOut[226]),
.io_out_227(dataOut[227]),
.io_out_228(dataOut[228]),
.io_out_229(dataOut[229]),
.io_out_230(dataOut[230]),
.io_out_231(dataOut[231]),
.io_out_232(dataOut[232]),
.io_out_233(dataOut[233]),
.io_out_234(dataOut[234]),
.io_out_235(dataOut[235]),
.io_out_236(dataOut[236]),
.io_out_237(dataOut[237]),
.io_out_238(dataOut[238]),
.io_out_239(dataOut[239]),
.io_out_240(dataOut[240]),
.io_out_241(dataOut[241]),
.io_out_242(dataOut[242]),
.io_out_243(dataOut[243]),
.io_out_244(dataOut[244]),
.io_out_245(dataOut[245]),
.io_out_246(dataOut[246]),
.io_out_247(dataOut[247]),
.io_out_248(dataOut[248]),
.io_out_249(dataOut[249]),
.io_out_250(dataOut[250]),
.io_out_251(dataOut[251]),
.io_out_252(dataOut[252]),
.io_out_253(dataOut[253]),
.io_out_254(dataOut[254]),
.io_out_255(dataOut[255]),
.io_out_256(dataOut[256]),
.io_out_257(dataOut[257]),
.io_out_258(dataOut[258]),
.io_out_259(dataOut[259]),
.io_out_260(dataOut[260]),
.io_out_261(dataOut[261]),
.io_out_262(dataOut[262]),
.io_out_263(dataOut[263]),
.io_out_264(dataOut[264]),
.io_out_265(dataOut[265]),
.io_out_266(dataOut[266]),
.io_out_267(dataOut[267]),
.io_out_268(dataOut[268]),
.io_out_269(dataOut[269]),
.io_out_270(dataOut[270]),
.io_out_271(dataOut[271]),
.io_out_272(dataOut[272]),
.io_out_273(dataOut[273]),
.io_out_274(dataOut[274]),
.io_out_275(dataOut[275]),
.io_out_276(dataOut[276]),
.io_out_277(dataOut[277]),
.io_out_278(dataOut[278]),
.io_out_279(dataOut[279]),
.io_out_280(dataOut[280]),
.io_out_281(dataOut[281]),
.io_out_282(dataOut[282]),
.io_out_283(dataOut[283]),
.io_out_284(dataOut[284]),
.io_out_285(dataOut[285]),
.io_out_286(dataOut[286]),
.io_out_287(dataOut[287]),
.io_out_288(dataOut[288]),
.io_out_289(dataOut[289]),
.io_out_290(dataOut[290]),
.io_out_291(dataOut[291]),
.io_out_292(dataOut[292]),
.io_out_293(dataOut[293]),
.io_out_294(dataOut[294]),
.io_out_295(dataOut[295]),
.io_out_296(dataOut[296]),
.io_out_297(dataOut[297]),
.io_out_298(dataOut[298]),
.io_out_299(dataOut[299]),
.io_out_300(dataOut[300]),
.io_out_301(dataOut[301]),
.io_out_302(dataOut[302]),
.io_out_303(dataOut[303]),
.io_out_304(dataOut[304]),
.io_out_305(dataOut[305]),
.io_out_306(dataOut[306]),
.io_out_307(dataOut[307]),
.io_out_308(dataOut[308]),
.io_out_309(dataOut[309]),
.io_out_310(dataOut[310]),
.io_out_311(dataOut[311]),
.io_out_312(dataOut[312]),
.io_out_313(dataOut[313]),
.io_out_314(dataOut[314]),
.io_out_315(dataOut[315]),
.io_out_316(dataOut[316]),
.io_out_317(dataOut[317]),
.io_out_318(dataOut[318]),
.io_out_319(dataOut[319]),
.io_out_320(dataOut[320]),
.io_out_321(dataOut[321]),
.io_out_322(dataOut[322]),
.io_out_323(dataOut[323]),
.io_out_324(dataOut[324]),
.io_out_325(dataOut[325]),
.io_out_326(dataOut[326]),
.io_out_327(dataOut[327]),
.io_out_328(dataOut[328]),
.io_out_329(dataOut[329]),
.io_out_330(dataOut[330]),
.io_out_331(dataOut[331]),
.io_out_332(dataOut[332]),
.io_out_333(dataOut[333]),
.io_out_334(dataOut[334]),
.io_out_335(dataOut[335]),
.io_out_336(dataOut[336]),
.io_out_337(dataOut[337]),
.io_out_338(dataOut[338]),
.io_out_339(dataOut[339]),
.io_out_340(dataOut[340]),
.io_out_341(dataOut[341]),
.io_out_342(dataOut[342]),
.io_out_343(dataOut[343]),
.io_out_344(dataOut[344]),
.io_out_345(dataOut[345]),
.io_out_346(dataOut[346]),
.io_out_347(dataOut[347]),
.io_out_348(dataOut[348]),
.io_out_349(dataOut[349]),
.io_out_350(dataOut[350]),
.io_out_351(dataOut[351]),
.io_out_352(dataOut[352]),
.io_out_353(dataOut[353]),
.io_out_354(dataOut[354]),
.io_out_355(dataOut[355]),
.io_out_356(dataOut[356]),
.io_out_357(dataOut[357]),
.io_out_358(dataOut[358]),
.io_out_359(dataOut[359]),
.io_out_360(dataOut[360]),
.io_out_361(dataOut[361]),
.io_out_362(dataOut[362]),
.io_out_363(dataOut[363]),
.io_out_364(dataOut[364]),
.io_out_365(dataOut[365]),
.io_out_366(dataOut[366]),
.io_out_367(dataOut[367]),
.io_out_368(dataOut[368]),
.io_out_369(dataOut[369]),
.io_out_370(dataOut[370]),
.io_out_371(dataOut[371]),
.io_out_372(dataOut[372]),
.io_out_373(dataOut[373]),
.io_out_374(dataOut[374]),
.io_out_375(dataOut[375]),
.io_out_376(dataOut[376]),
.io_out_377(dataOut[377]),
.io_out_378(dataOut[378]),
.io_out_379(dataOut[379]),
.io_out_380(dataOut[380]),
.io_out_381(dataOut[381]),
.io_out_382(dataOut[382]),
.io_out_383(dataOut[383]),
.io_out_384(dataOut[384]),
.io_out_385(dataOut[385]),
.io_out_386(dataOut[386]),
.io_out_387(dataOut[387]),
.io_out_388(dataOut[388]),
.io_out_389(dataOut[389]),
.io_out_390(dataOut[390]),
.io_out_391(dataOut[391]),
.io_out_392(dataOut[392]),
.io_out_393(dataOut[393]),
.io_out_394(dataOut[394]),
.io_out_395(dataOut[395]),
.io_out_396(dataOut[396]),
.io_out_397(dataOut[397]),
.io_out_398(dataOut[398]),
.io_out_399(dataOut[399]),
.io_out_400(dataOut[400]),
.io_out_401(dataOut[401]),
.io_out_402(dataOut[402]),
.io_out_403(dataOut[403]),
.io_out_404(dataOut[404]),
.io_out_405(dataOut[405]),
.io_out_406(dataOut[406]),
.io_out_407(dataOut[407]),
.io_out_408(dataOut[408]),
.io_out_409(dataOut[409]),
.io_out_410(dataOut[410]),
.io_out_411(dataOut[411]),
.io_out_412(dataOut[412]),
.io_out_413(dataOut[413]),
.io_out_414(dataOut[414]),
.io_out_415(dataOut[415]),
.io_out_416(dataOut[416]),
.io_out_417(dataOut[417]),
.io_out_418(dataOut[418]),
.io_out_419(dataOut[419]),
.io_out_420(dataOut[420]),
.io_out_421(dataOut[421]),
.io_out_422(dataOut[422]),
.io_out_423(dataOut[423]),
.io_out_424(dataOut[424]),
.io_out_425(dataOut[425]),
.io_out_426(dataOut[426]),
.io_out_427(dataOut[427]),
.io_out_428(dataOut[428]),
.io_out_429(dataOut[429]),
.io_out_430(dataOut[430]),
.io_out_431(dataOut[431]),
.io_out_432(dataOut[432]),
.io_out_433(dataOut[433]),
.io_out_434(dataOut[434]),
.io_out_435(dataOut[435]),
.io_out_436(dataOut[436]),
.io_out_437(dataOut[437]),
.io_out_438(dataOut[438]),
.io_out_439(dataOut[439]),
.io_out_440(dataOut[440]),
.io_out_441(dataOut[441]),
.io_out_442(dataOut[442]),
.io_out_443(dataOut[443]),
.io_out_444(dataOut[444]),
.io_out_445(dataOut[445]),
.io_out_446(dataOut[446]),
.io_out_447(dataOut[447]),
.io_out_448(dataOut[448]),
.io_out_449(dataOut[449]),
.io_out_450(dataOut[450]),
.io_out_451(dataOut[451]),
.io_out_452(dataOut[452]),
.io_out_453(dataOut[453]),
.io_out_454(dataOut[454]),
.io_out_455(dataOut[455]),
.io_out_456(dataOut[456]),
.io_out_457(dataOut[457]),
.io_out_458(dataOut[458]),
.io_out_459(dataOut[459]),
.io_out_460(dataOut[460]),
.io_out_461(dataOut[461]),
.io_out_462(dataOut[462]),
.io_out_463(dataOut[463]),
.io_out_464(dataOut[464]),
.io_out_465(dataOut[465]),
.io_out_466(dataOut[466]),
.io_out_467(dataOut[467]),
.io_out_468(dataOut[468]),
.io_out_469(dataOut[469]),
.io_out_470(dataOut[470]),
.io_out_471(dataOut[471]),
.io_out_472(dataOut[472]),
.io_out_473(dataOut[473]),
.io_out_474(dataOut[474]),
.io_out_475(dataOut[475]),
.io_out_476(dataOut[476]),
.io_out_477(dataOut[477]),
.io_out_478(dataOut[478]),
.io_out_479(dataOut[479]),
.io_out_480(dataOut[480]),
.io_out_481(dataOut[481]),
.io_out_482(dataOut[482]),
.io_out_483(dataOut[483]),
.io_out_484(dataOut[484]),
.io_out_485(dataOut[485]),
.io_out_486(dataOut[486]),
.io_out_487(dataOut[487]),
.io_out_488(dataOut[488]),
.io_out_489(dataOut[489]),
.io_out_490(dataOut[490]),
.io_out_491(dataOut[491]),
.io_out_492(dataOut[492]),
.io_out_493(dataOut[493]),
.io_out_494(dataOut[494]),
.io_out_495(dataOut[495]),
.io_out_496(dataOut[496]),
.io_out_497(dataOut[497]),
.io_out_498(dataOut[498]),
.io_out_499(dataOut[499]),
.io_out_500(dataOut[500]),
.io_out_501(dataOut[501]),
.io_out_502(dataOut[502]),
.io_out_503(dataOut[503]),
.io_out_504(dataOut[504]),
.io_out_505(dataOut[505]),
.io_out_506(dataOut[506]),
.io_out_507(dataOut[507]),
.io_out_508(dataOut[508]),
.io_out_509(dataOut[509]),
.io_out_510(dataOut[510]),
.io_out_511(dataOut[511]),
.io_out_512(dataOut[512]),
.io_out_513(dataOut[513]),
.io_out_514(dataOut[514]),
.io_out_515(dataOut[515]),
.io_out_516(dataOut[516]),
.io_out_517(dataOut[517]),
.io_out_518(dataOut[518]),
.io_out_519(dataOut[519]),
.io_out_520(dataOut[520]),
.io_out_521(dataOut[521]),
.io_out_522(dataOut[522]),
.io_out_523(dataOut[523]),
.io_out_524(dataOut[524]),
.io_out_525(dataOut[525]),
.io_out_526(dataOut[526]),
.io_out_527(dataOut[527]),
.io_out_528(dataOut[528]),
.io_out_529(dataOut[529]),
.io_out_530(dataOut[530]),
.io_out_531(dataOut[531]),
.io_out_532(dataOut[532]),
.io_out_533(dataOut[533]),
.io_out_534(dataOut[534]),
.io_out_535(dataOut[535]),
.io_out_536(dataOut[536]),
.io_out_537(dataOut[537]),
.io_out_538(dataOut[538]),
.io_out_539(dataOut[539]),
.io_out_540(dataOut[540]),
.io_out_541(dataOut[541]),
.io_out_542(dataOut[542]),
.io_out_543(dataOut[543]),
.io_out_544(dataOut[544]),
.io_out_545(dataOut[545]),
.io_out_546(dataOut[546]),
.io_out_547(dataOut[547]),
.io_out_548(dataOut[548]),
.io_out_549(dataOut[549]),
.io_out_550(dataOut[550]),
.io_out_551(dataOut[551]),
.io_out_552(dataOut[552]),
.io_out_553(dataOut[553]),
.io_out_554(dataOut[554]),
.io_out_555(dataOut[555]),
.io_out_556(dataOut[556]),
.io_out_557(dataOut[557]),
.io_out_558(dataOut[558]),
.io_out_559(dataOut[559]),
.io_out_560(dataOut[560]),
.io_out_561(dataOut[561]),
.io_out_562(dataOut[562]),
.io_out_563(dataOut[563]),
.io_out_564(dataOut[564]),
.io_out_565(dataOut[565]),
.io_out_566(dataOut[566]),
.io_out_567(dataOut[567]),
.io_out_568(dataOut[568]),
.io_out_569(dataOut[569]),
.io_out_570(dataOut[570]),
.io_out_571(dataOut[571]),
.io_out_572(dataOut[572]),
.io_out_573(dataOut[573]),
.io_out_574(dataOut[574]),
.io_out_575(dataOut[575]),
.io_out_576(dataOut[576]),
.io_out_577(dataOut[577]),
.io_out_578(dataOut[578]),
.io_out_579(dataOut[579]),
.io_out_580(dataOut[580]),
.io_out_581(dataOut[581]),
.io_out_582(dataOut[582]),
.io_out_583(dataOut[583]),
.io_out_584(dataOut[584]),
.io_out_585(dataOut[585]),
.io_out_586(dataOut[586]),
.io_out_587(dataOut[587]),
.io_out_588(dataOut[588]),
.io_out_589(dataOut[589]),
.io_out_590(dataOut[590]),
.io_out_591(dataOut[591]),
.io_out_592(dataOut[592]),
.io_out_593(dataOut[593]),
.io_out_594(dataOut[594]),
.io_out_595(dataOut[595]),
.io_out_596(dataOut[596]),
.io_out_597(dataOut[597]),
.io_out_598(dataOut[598]),
.io_out_599(dataOut[599]),
.io_out_600(dataOut[600]),
.io_out_601(dataOut[601]),
.io_out_602(dataOut[602]),
.io_out_603(dataOut[603]),
.io_out_604(dataOut[604]),
.io_out_605(dataOut[605]),
.io_out_606(dataOut[606]),
.io_out_607(dataOut[607]),
.io_out_608(dataOut[608]),
.io_out_609(dataOut[609]),
.io_out_610(dataOut[610]),
.io_out_611(dataOut[611]),
.io_out_612(dataOut[612]),
.io_out_613(dataOut[613]),
.io_out_614(dataOut[614]),
.io_out_615(dataOut[615]),
.io_out_616(dataOut[616]),
.io_out_617(dataOut[617]),
.io_out_618(dataOut[618]),
.io_out_619(dataOut[619]),
.io_out_620(dataOut[620]),
.io_out_621(dataOut[621]),
.io_out_622(dataOut[622]),
.io_out_623(dataOut[623]),
.io_out_624(dataOut[624]),
.io_out_625(dataOut[625]),
.io_out_626(dataOut[626]),
.io_out_627(dataOut[627]),
.io_out_628(dataOut[628]),
.io_out_629(dataOut[629]),
.io_out_630(dataOut[630]),
.io_out_631(dataOut[631]),
.io_out_632(dataOut[632]),
.io_out_633(dataOut[633]),
.io_out_634(dataOut[634]),
.io_out_635(dataOut[635]),
.io_out_636(dataOut[636]),
.io_out_637(dataOut[637]),
.io_out_638(dataOut[638]),
.io_out_639(dataOut[639]),
.io_out_640(dataOut[640]),
.io_out_641(dataOut[641]),
.io_out_642(dataOut[642]),
.io_out_643(dataOut[643]),
.io_out_644(dataOut[644]),
.io_out_645(dataOut[645]),
.io_out_646(dataOut[646]),
.io_out_647(dataOut[647]),
.io_out_648(dataOut[648]),
.io_out_649(dataOut[649]),
.io_out_650(dataOut[650]),
.io_out_651(dataOut[651]),
.io_out_652(dataOut[652]),
.io_out_653(dataOut[653]),
.io_out_654(dataOut[654]),
.io_out_655(dataOut[655]),
.io_out_656(dataOut[656]),
.io_out_657(dataOut[657]),
.io_out_658(dataOut[658]),
.io_out_659(dataOut[659]),
.io_out_660(dataOut[660]),
.io_out_661(dataOut[661]),
.io_out_662(dataOut[662]),
.io_out_663(dataOut[663]),
.io_out_664(dataOut[664]),
.io_out_665(dataOut[665]),
.io_out_666(dataOut[666]),
.io_out_667(dataOut[667]),
.io_out_668(dataOut[668]),
.io_out_669(dataOut[669]),
.io_out_670(dataOut[670]),
.io_out_671(dataOut[671]),
.io_out_672(dataOut[672]),
.io_out_673(dataOut[673]),
.io_out_674(dataOut[674]),
.io_out_675(dataOut[675]),
.io_out_676(dataOut[676]),
.io_out_677(dataOut[677]),
.io_out_678(dataOut[678]),
.io_out_679(dataOut[679]),
.io_out_680(dataOut[680]),
.io_out_681(dataOut[681]),
.io_out_682(dataOut[682]),
.io_out_683(dataOut[683]),
.io_out_684(dataOut[684]),
.io_out_685(dataOut[685]),
.io_out_686(dataOut[686]),
.io_out_687(dataOut[687]),
.io_out_688(dataOut[688]),
.io_out_689(dataOut[689]),
.io_out_690(dataOut[690]),
.io_out_691(dataOut[691]),
.io_out_692(dataOut[692]),
.io_out_693(dataOut[693]),
.io_out_694(dataOut[694]),
.io_out_695(dataOut[695]),
.io_out_696(dataOut[696]),
.io_out_697(dataOut[697]),
.io_out_698(dataOut[698]),
.io_out_699(dataOut[699]),
.io_out_700(dataOut[700]),
.io_out_701(dataOut[701]),
.io_out_702(dataOut[702]),
.io_out_703(dataOut[703]),
.io_out_704(dataOut[704]),
.io_out_705(dataOut[705]),
.io_out_706(dataOut[706]),
.io_out_707(dataOut[707]),
.io_out_708(dataOut[708]),
.io_out_709(dataOut[709]),
.io_out_710(dataOut[710]),
.io_out_711(dataOut[711]),
.io_out_712(dataOut[712]),
.io_out_713(dataOut[713]),
.io_out_714(dataOut[714]),
.io_out_715(dataOut[715]),
.io_out_716(dataOut[716]),
.io_out_717(dataOut[717]),
.io_out_718(dataOut[718]),
.io_out_719(dataOut[719]),
.io_out_720(dataOut[720]),
.io_out_721(dataOut[721]),
.io_out_722(dataOut[722]),
.io_out_723(dataOut[723]),
.io_out_724(dataOut[724]),
.io_out_725(dataOut[725]),
.io_out_726(dataOut[726]),
.io_out_727(dataOut[727]),
.io_out_728(dataOut[728]),
.io_out_729(dataOut[729]),
.io_out_730(dataOut[730]),
.io_out_731(dataOut[731]),
.io_out_732(dataOut[732]),
.io_out_733(dataOut[733]),
.io_out_734(dataOut[734]),
.io_out_735(dataOut[735]),
.io_out_736(dataOut[736]),
.io_out_737(dataOut[737]),
.io_out_738(dataOut[738]),
.io_out_739(dataOut[739]),
.io_out_740(dataOut[740]),
.io_out_741(dataOut[741]),
.io_out_742(dataOut[742]),
.io_out_743(dataOut[743]),
.io_out_744(dataOut[744]),
.io_out_745(dataOut[745]),
.io_out_746(dataOut[746]),
.io_out_747(dataOut[747]),
.io_out_748(dataOut[748]),
.io_out_749(dataOut[749]),
.io_out_750(dataOut[750]),
.io_out_751(dataOut[751]),
.io_out_752(dataOut[752]),
.io_out_753(dataOut[753]),
.io_out_754(dataOut[754]),
.io_out_755(dataOut[755]),
.io_out_756(dataOut[756]),
.io_out_757(dataOut[757]),
.io_out_758(dataOut[758]),
.io_out_759(dataOut[759]),
.io_out_760(dataOut[760]),
.io_out_761(dataOut[761]),
.io_out_762(dataOut[762]),
.io_out_763(dataOut[763]),
.io_out_764(dataOut[764]),
.io_out_765(dataOut[765]),
.io_out_766(dataOut[766]),
.io_out_767(dataOut[767]),
.io_out_768(dataOut[768]),
.io_out_769(dataOut[769]),
.io_out_770(dataOut[770]),
.io_out_771(dataOut[771]),
.io_out_772(dataOut[772]),
.io_out_773(dataOut[773]),
.io_out_774(dataOut[774]),
.io_out_775(dataOut[775]),
.io_out_776(dataOut[776]),
.io_out_777(dataOut[777]),
.io_out_778(dataOut[778]),
.io_out_779(dataOut[779]),
.io_out_780(dataOut[780]),
.io_out_781(dataOut[781]),
.io_out_782(dataOut[782]),
.io_out_783(dataOut[783]),
.io_out_784(dataOut[784]),
.io_out_785(dataOut[785]),
.io_out_786(dataOut[786]),
.io_out_787(dataOut[787]),
.io_out_788(dataOut[788]),
.io_out_789(dataOut[789]),
.io_out_790(dataOut[790]),
.io_out_791(dataOut[791]),
.io_out_792(dataOut[792]),
.io_out_793(dataOut[793]),
.io_out_794(dataOut[794]),
.io_out_795(dataOut[795]),
.io_out_796(dataOut[796]),
.io_out_797(dataOut[797]),
.io_out_798(dataOut[798]),
.io_out_799(dataOut[799]),
.io_out_800(dataOut[800]),
.io_out_801(dataOut[801]),
.io_out_802(dataOut[802]),
.io_out_803(dataOut[803]),
.io_out_804(dataOut[804]),
.io_out_805(dataOut[805]),
.io_out_806(dataOut[806]),
.io_out_807(dataOut[807]),
.io_out_808(dataOut[808]),
.io_out_809(dataOut[809]),
.io_out_810(dataOut[810]),
.io_out_811(dataOut[811]),
.io_out_812(dataOut[812]),
.io_out_813(dataOut[813]),
.io_out_814(dataOut[814]),
.io_out_815(dataOut[815]),
.io_out_816(dataOut[816]),
.io_out_817(dataOut[817]),
.io_out_818(dataOut[818]),
.io_out_819(dataOut[819]),
.io_out_820(dataOut[820]),
.io_out_821(dataOut[821]),
.io_out_822(dataOut[822]),
.io_out_823(dataOut[823]),
.io_out_824(dataOut[824]),
.io_out_825(dataOut[825]),
.io_out_826(dataOut[826]),
.io_out_827(dataOut[827]),
.io_out_828(dataOut[828]),
.io_out_829(dataOut[829]),
.io_out_830(dataOut[830]),
.io_out_831(dataOut[831]),
.io_out_832(dataOut[832]),
.io_out_833(dataOut[833]),
.io_out_834(dataOut[834]),
.io_out_835(dataOut[835]),
.io_out_836(dataOut[836]),
.io_out_837(dataOut[837]),
.io_out_838(dataOut[838]),
.io_out_839(dataOut[839]),
.io_out_840(dataOut[840]),
.io_out_841(dataOut[841]),
.io_out_842(dataOut[842]),
.io_out_843(dataOut[843]),
.io_out_844(dataOut[844]),
.io_out_845(dataOut[845]),
.io_out_846(dataOut[846]),
.io_out_847(dataOut[847]),
.io_out_848(dataOut[848]),
.io_out_849(dataOut[849]),
.io_out_850(dataOut[850]),
.io_out_851(dataOut[851]),
.io_out_852(dataOut[852]),
.io_out_853(dataOut[853]),
.io_out_854(dataOut[854]),
.io_out_855(dataOut[855]),
.io_out_856(dataOut[856]),
.io_out_857(dataOut[857]),
.io_out_858(dataOut[858]),
.io_out_859(dataOut[859]),
.io_out_860(dataOut[860]),
.io_out_861(dataOut[861]),
.io_out_862(dataOut[862]),
.io_out_863(dataOut[863]),
.io_out_864(dataOut[864]),
.io_out_865(dataOut[865]),
.io_out_866(dataOut[866]),
.io_out_867(dataOut[867]),
.io_out_868(dataOut[868]),
.io_out_869(dataOut[869]),
.io_out_870(dataOut[870]),
.io_out_871(dataOut[871]),
.io_out_872(dataOut[872]),
.io_out_873(dataOut[873]),
.io_out_874(dataOut[874]),
.io_out_875(dataOut[875]),
.io_out_876(dataOut[876]),
.io_out_877(dataOut[877]),
.io_out_878(dataOut[878]),
.io_out_879(dataOut[879]),
.io_out_880(dataOut[880]),
.io_out_881(dataOut[881]),
.io_out_882(dataOut[882]),
.io_out_883(dataOut[883]),
.io_out_884(dataOut[884]),
.io_out_885(dataOut[885]),
.io_out_886(dataOut[886]),
.io_out_887(dataOut[887]),
.io_out_888(dataOut[888]),
.io_out_889(dataOut[889]),
.io_out_890(dataOut[890]),
.io_out_891(dataOut[891]),
.io_out_892(dataOut[892]),
.io_out_893(dataOut[893]),
.io_out_894(dataOut[894]),
.io_out_895(dataOut[895]),
.io_out_896(dataOut[896]),
.io_out_897(dataOut[897]),
.io_out_898(dataOut[898]),
.io_out_899(dataOut[899]),
.io_out_900(dataOut[900]),
.io_out_901(dataOut[901]),
.io_out_902(dataOut[902]),
.io_out_903(dataOut[903]),
.io_out_904(dataOut[904]),
.io_out_905(dataOut[905]),
.io_out_906(dataOut[906]),
.io_out_907(dataOut[907]),
.io_out_908(dataOut[908]),
.io_out_909(dataOut[909]),
.io_out_910(dataOut[910]),
.io_out_911(dataOut[911]),
.io_out_912(dataOut[912]),
.io_out_913(dataOut[913]),
.io_out_914(dataOut[914]),
.io_out_915(dataOut[915]),
.io_out_916(dataOut[916]),
.io_out_917(dataOut[917]),
.io_out_918(dataOut[918]),
.io_out_919(dataOut[919]),
.io_out_920(dataOut[920]),
.io_out_921(dataOut[921]),
.io_out_922(dataOut[922]),
.io_out_923(dataOut[923]),
.io_out_924(dataOut[924]),
.io_out_925(dataOut[925]),
.io_out_926(dataOut[926]),
.io_out_927(dataOut[927]),
.io_out_928(dataOut[928]),
.io_out_929(dataOut[929]),
.io_out_930(dataOut[930]),
.io_out_931(dataOut[931]),
.io_out_932(dataOut[932]),
.io_out_933(dataOut[933]),
.io_out_934(dataOut[934]),
.io_out_935(dataOut[935]),
.io_out_936(dataOut[936]),
.io_out_937(dataOut[937]),
.io_out_938(dataOut[938]),
.io_out_939(dataOut[939]),
.io_out_940(dataOut[940]),
.io_out_941(dataOut[941]),
.io_out_942(dataOut[942]),
.io_out_943(dataOut[943]),
.io_out_944(dataOut[944]),
.io_out_945(dataOut[945]),
.io_out_946(dataOut[946]),
.io_out_947(dataOut[947]),
.io_out_948(dataOut[948]),
.io_out_949(dataOut[949]),
.io_out_950(dataOut[950]),
.io_out_951(dataOut[951]),
.io_out_952(dataOut[952]),
.io_out_953(dataOut[953]),
.io_out_954(dataOut[954]),
.io_out_955(dataOut[955]),
.io_out_956(dataOut[956]),
.io_out_957(dataOut[957]),
.io_out_958(dataOut[958]),
.io_out_959(dataOut[959]),
.io_out_960(dataOut[960]),
.io_out_961(dataOut[961]),
.io_out_962(dataOut[962]),
.io_out_963(dataOut[963]),
.io_out_964(dataOut[964]),
.io_out_965(dataOut[965]),
.io_out_966(dataOut[966]),
.io_out_967(dataOut[967]),
.io_out_968(dataOut[968]),
.io_out_969(dataOut[969]),
.io_out_970(dataOut[970]),
.io_out_971(dataOut[971]),
.io_out_972(dataOut[972]),
.io_out_973(dataOut[973]),
.io_out_974(dataOut[974]),
.io_out_975(dataOut[975]),
.io_out_976(dataOut[976]),
.io_out_977(dataOut[977]),
.io_out_978(dataOut[978]),
.io_out_979(dataOut[979]),
.io_out_980(dataOut[980]),
.io_out_981(dataOut[981]),
.io_out_982(dataOut[982]),
.io_out_983(dataOut[983]),
.io_out_984(dataOut[984]),
.io_out_985(dataOut[985]),
.io_out_986(dataOut[986]),
.io_out_987(dataOut[987]),
.io_out_988(dataOut[988]),
.io_out_989(dataOut[989]),
.io_out_990(dataOut[990]),
.io_out_991(dataOut[991]),
.io_out_992(dataOut[992]),
.io_out_993(dataOut[993]),
.io_out_994(dataOut[994]),
.io_out_995(dataOut[995]),
.io_out_996(dataOut[996]),
.io_out_997(dataOut[997]),
.io_out_998(dataOut[998]),
.io_out_999(dataOut[999]),
.io_out_1000(dataOut[1000]),
.io_out_1001(dataOut[1001]),
.io_out_1002(dataOut[1002]),
.io_out_1003(dataOut[1003]),
.io_out_1004(dataOut[1004]),
.io_out_1005(dataOut[1005]),
.io_out_1006(dataOut[1006]),
.io_out_1007(dataOut[1007]),
.io_out_1008(dataOut[1008]),
.io_out_1009(dataOut[1009]),
.io_out_1010(dataOut[1010]),
.io_out_1011(dataOut[1011]),
.io_out_1012(dataOut[1012]),
.io_out_1013(dataOut[1013]),
.io_out_1014(dataOut[1014]),
.io_out_1015(dataOut[1015]),
.io_out_1016(dataOut[1016]),
.io_out_1017(dataOut[1017]),
.io_out_1018(dataOut[1018]),
.io_out_1019(dataOut[1019]),
.io_out_1020(dataOut[1020]),
.io_out_1021(dataOut[1021]),
.io_out_1022(dataOut[1022]),
.io_out_1023(dataOut[1023]),
.io_out_1024(dataOut[1024]),
.io_out_1025(dataOut[1025]),
.io_out_1026(dataOut[1026]),
.io_out_1027(dataOut[1027]),
.io_out_1028(dataOut[1028]),
.io_out_1029(dataOut[1029]),
.io_out_1030(dataOut[1030]),
.io_out_1031(dataOut[1031]),
.io_out_1032(dataOut[1032]),
.io_out_1033(dataOut[1033]),
.io_out_1034(dataOut[1034]),
.io_out_1035(dataOut[1035]),
.io_out_1036(dataOut[1036]),
.io_out_1037(dataOut[1037]),
.io_out_1038(dataOut[1038]),
.io_out_1039(dataOut[1039]),
.io_out_1040(dataOut[1040]),
.io_out_1041(dataOut[1041]),
.io_out_1042(dataOut[1042]),
.io_out_1043(dataOut[1043]),
.io_out_1044(dataOut[1044]),
.io_out_1045(dataOut[1045]),
.io_out_1046(dataOut[1046]),
.io_out_1047(dataOut[1047]),
.io_out_1048(dataOut[1048]),
.io_out_1049(dataOut[1049]),
.io_out_1050(dataOut[1050]),
.io_out_1051(dataOut[1051]),
.io_out_1052(dataOut[1052]),
.io_out_1053(dataOut[1053]),
.io_out_1054(dataOut[1054]),
.io_out_1055(dataOut[1055]),
.io_out_1056(dataOut[1056]),
.io_out_1057(dataOut[1057]),
.io_out_1058(dataOut[1058]),
.io_out_1059(dataOut[1059]),
.io_out_1060(dataOut[1060]),
.io_out_1061(dataOut[1061]),
.io_out_1062(dataOut[1062]),
.io_out_1063(dataOut[1063]),
.io_out_1064(dataOut[1064]),
.io_out_1065(dataOut[1065]),
.io_out_1066(dataOut[1066]),
.io_out_1067(dataOut[1067]),
.io_out_1068(dataOut[1068]),
.io_out_1069(dataOut[1069]),
.io_out_1070(dataOut[1070]),
.io_out_1071(dataOut[1071]),
.io_out_1072(dataOut[1072]),
.io_out_1073(dataOut[1073]),
.io_out_1074(dataOut[1074]),
.io_out_1075(dataOut[1075]),
.io_out_1076(dataOut[1076]),
.io_out_1077(dataOut[1077]),
.io_out_1078(dataOut[1078]),
.io_out_1079(dataOut[1079]),
.io_out_1080(dataOut[1080]),
.io_out_1081(dataOut[1081]),
.io_out_1082(dataOut[1082]),
.io_out_1083(dataOut[1083]),
.io_out_1084(dataOut[1084]),
.io_out_1085(dataOut[1085]),
.io_out_1086(dataOut[1086]),
.io_out_1087(dataOut[1087]),
.io_out_1088(dataOut[1088]),
.io_out_1089(dataOut[1089]),
.io_out_1090(dataOut[1090]),
.io_out_1091(dataOut[1091]),
.io_out_1092(dataOut[1092]),
.io_out_1093(dataOut[1093]),
.io_out_1094(dataOut[1094]),
.io_out_1095(dataOut[1095]),
.io_out_1096(dataOut[1096]),
.io_out_1097(dataOut[1097]),
.io_out_1098(dataOut[1098]),
.io_out_1099(dataOut[1099]),
.io_out_1100(dataOut[1100]),
.io_out_1101(dataOut[1101]),
.io_out_1102(dataOut[1102]),
.io_out_1103(dataOut[1103]),
.io_out_1104(dataOut[1104]),
.io_out_1105(dataOut[1105]),
.io_out_1106(dataOut[1106]),
.io_out_1107(dataOut[1107]),
.io_out_1108(dataOut[1108]),
.io_out_1109(dataOut[1109]),
.io_out_1110(dataOut[1110]),
.io_out_1111(dataOut[1111]),
.io_out_1112(dataOut[1112]),
.io_out_1113(dataOut[1113]),
.io_out_1114(dataOut[1114]),
.io_out_1115(dataOut[1115]),
.io_out_1116(dataOut[1116]),
.io_out_1117(dataOut[1117]),
.io_out_1118(dataOut[1118]),
.io_out_1119(dataOut[1119]),
.io_out_1120(dataOut[1120]),
.io_out_1121(dataOut[1121]),
.io_out_1122(dataOut[1122]),
.io_out_1123(dataOut[1123]),
.io_out_1124(dataOut[1124]),
.io_out_1125(dataOut[1125]),
.io_out_1126(dataOut[1126]),
.io_out_1127(dataOut[1127]),
.io_out_1128(dataOut[1128]),
.io_out_1129(dataOut[1129]),
.io_out_1130(dataOut[1130]),
.io_out_1131(dataOut[1131]),
.io_out_1132(dataOut[1132]),
.io_out_1133(dataOut[1133]),
.io_out_1134(dataOut[1134]),
.io_out_1135(dataOut[1135]),
.io_out_1136(dataOut[1136]),
.io_out_1137(dataOut[1137]),
.io_out_1138(dataOut[1138]),
.io_out_1139(dataOut[1139]),
.io_out_1140(dataOut[1140]),
.io_out_1141(dataOut[1141]),
.io_out_1142(dataOut[1142]),
.io_out_1143(dataOut[1143]),
.io_out_1144(dataOut[1144]),
.io_out_1145(dataOut[1145]),
.io_out_1146(dataOut[1146]),
.io_out_1147(dataOut[1147]),
.io_out_1148(dataOut[1148]),
.io_out_1149(dataOut[1149]),
.io_out_1150(dataOut[1150]),
.io_out_1151(dataOut[1151]),
.io_out_1152(dataOut[1152]),
.io_out_1153(dataOut[1153]),
.io_out_1154(dataOut[1154]),
.io_out_1155(dataOut[1155]),
.io_out_1156(dataOut[1156]),
.io_out_1157(dataOut[1157]),
.io_out_1158(dataOut[1158]),
.io_out_1159(dataOut[1159]),
.io_out_1160(dataOut[1160]),
.io_out_1161(dataOut[1161]),
.io_out_1162(dataOut[1162]),
.io_out_1163(dataOut[1163]),
.io_out_1164(dataOut[1164]),
.io_out_1165(dataOut[1165]),
.io_out_1166(dataOut[1166]),
.io_out_1167(dataOut[1167]),
.io_out_1168(dataOut[1168]),
.io_out_1169(dataOut[1169]),
.io_out_1170(dataOut[1170]),
.io_out_1171(dataOut[1171]),
.io_out_1172(dataOut[1172]),
.io_out_1173(dataOut[1173]),
.io_out_1174(dataOut[1174]),
.io_out_1175(dataOut[1175]),
.io_out_1176(dataOut[1176]),
.io_out_1177(dataOut[1177]),
.io_out_1178(dataOut[1178]),
.io_out_1179(dataOut[1179]),
.io_out_1180(dataOut[1180]),
.io_out_1181(dataOut[1181]),
.io_out_1182(dataOut[1182]),
.io_out_1183(dataOut[1183]),
.io_out_1184(dataOut[1184]),
.io_out_1185(dataOut[1185]),
.io_out_1186(dataOut[1186]),
.io_out_1187(dataOut[1187]),
.io_out_1188(dataOut[1188]),
.io_out_1189(dataOut[1189]),
.io_out_1190(dataOut[1190]),
.io_out_1191(dataOut[1191]),
.io_out_1192(dataOut[1192]),
.io_out_1193(dataOut[1193]),
.io_out_1194(dataOut[1194]),
.io_out_1195(dataOut[1195]),
.io_out_1196(dataOut[1196]),
.io_out_1197(dataOut[1197]),
.io_out_1198(dataOut[1198]),
.io_out_1199(dataOut[1199]),
.io_out_1200(dataOut[1200]),
.io_out_1201(dataOut[1201]),
.io_out_1202(dataOut[1202]),
.io_out_1203(dataOut[1203]),
.io_out_1204(dataOut[1204]),
.io_out_1205(dataOut[1205]),
.io_out_1206(dataOut[1206]),
.io_out_1207(dataOut[1207]),
.io_out_1208(dataOut[1208]),
.io_out_1209(dataOut[1209]),
.io_out_1210(dataOut[1210]),
.io_out_1211(dataOut[1211]),
.io_out_1212(dataOut[1212]),
.io_out_1213(dataOut[1213]),
.io_out_1214(dataOut[1214]),
.io_out_1215(dataOut[1215]),
.io_out_1216(dataOut[1216]),
.io_out_1217(dataOut[1217]),
.io_out_1218(dataOut[1218]),
.io_out_1219(dataOut[1219]),
.io_out_1220(dataOut[1220]),
.io_out_1221(dataOut[1221]),
.io_out_1222(dataOut[1222]),
.io_out_1223(dataOut[1223]),
.io_out_1224(dataOut[1224]),
.io_out_1225(dataOut[1225]),
.io_out_1226(dataOut[1226]),
.io_out_1227(dataOut[1227]),
.io_out_1228(dataOut[1228]),
.io_out_1229(dataOut[1229]),
.io_out_1230(dataOut[1230]),
.io_out_1231(dataOut[1231]),
.io_out_1232(dataOut[1232]),
.io_out_1233(dataOut[1233]),
.io_out_1234(dataOut[1234]),
.io_out_1235(dataOut[1235]),
.io_out_1236(dataOut[1236]),
.io_out_1237(dataOut[1237]),
.io_out_1238(dataOut[1238]),
.io_out_1239(dataOut[1239]),
.io_out_1240(dataOut[1240]),
.io_out_1241(dataOut[1241]),
.io_out_1242(dataOut[1242]),
.io_out_1243(dataOut[1243]),
.io_out_1244(dataOut[1244]),
.io_out_1245(dataOut[1245]),
.io_out_1246(dataOut[1246]),
.io_out_1247(dataOut[1247]),
.io_out_1248(dataOut[1248]),
.io_out_1249(dataOut[1249]),
.io_out_1250(dataOut[1250]),
.io_out_1251(dataOut[1251]),
.io_out_1252(dataOut[1252]),
.io_out_1253(dataOut[1253]),
.io_out_1254(dataOut[1254]),
.io_out_1255(dataOut[1255]),
.io_out_1256(dataOut[1256]),
.io_out_1257(dataOut[1257]),
.io_out_1258(dataOut[1258]),
.io_out_1259(dataOut[1259]),
.io_out_1260(dataOut[1260]),
.io_out_1261(dataOut[1261]),
.io_out_1262(dataOut[1262]),
.io_out_1263(dataOut[1263]),
.io_out_1264(dataOut[1264]),
.io_out_1265(dataOut[1265]),
.io_out_1266(dataOut[1266]),
.io_out_1267(dataOut[1267]),
.io_out_1268(dataOut[1268]),
.io_out_1269(dataOut[1269]),
.io_out_1270(dataOut[1270]),
.io_out_1271(dataOut[1271]),
.io_out_1272(dataOut[1272]),
.io_out_1273(dataOut[1273]),
.io_out_1274(dataOut[1274]),
.io_out_1275(dataOut[1275]),
.io_out_1276(dataOut[1276]),
.io_out_1277(dataOut[1277]),
.io_out_1278(dataOut[1278]),
.io_out_1279(dataOut[1279]),
.io_out_1280(dataOut[1280]),
.io_out_1281(dataOut[1281]),
.io_out_1282(dataOut[1282]),
.io_out_1283(dataOut[1283]),
.io_out_1284(dataOut[1284]),
.io_out_1285(dataOut[1285]),
.io_out_1286(dataOut[1286]),
.io_out_1287(dataOut[1287]),
.io_out_1288(dataOut[1288]),
.io_out_1289(dataOut[1289]),
.io_out_1290(dataOut[1290]),
.io_out_1291(dataOut[1291]),
.io_out_1292(dataOut[1292]),
.io_out_1293(dataOut[1293]),
.io_out_1294(dataOut[1294]),
.io_out_1295(dataOut[1295]),
.io_out_1296(dataOut[1296]),
.io_out_1297(dataOut[1297]),
.io_out_1298(dataOut[1298]),
.io_out_1299(dataOut[1299]),
.io_out_1300(dataOut[1300]),
.io_out_1301(dataOut[1301]),
.io_out_1302(dataOut[1302]),
.io_out_1303(dataOut[1303]),
.io_out_1304(dataOut[1304]),
.io_out_1305(dataOut[1305]),
.io_out_1306(dataOut[1306]),
.io_out_1307(dataOut[1307]),
.io_out_1308(dataOut[1308]),
.io_out_1309(dataOut[1309]),
.io_out_1310(dataOut[1310]),
.io_out_1311(dataOut[1311]),
.io_out_1312(dataOut[1312]),
.io_out_1313(dataOut[1313]),
.io_out_1314(dataOut[1314]),
.io_out_1315(dataOut[1315]),
.io_out_1316(dataOut[1316]),
.io_out_1317(dataOut[1317]),
.io_out_1318(dataOut[1318]),
.io_out_1319(dataOut[1319]),
.io_out_1320(dataOut[1320]),
.io_out_1321(dataOut[1321]),
.io_out_1322(dataOut[1322]),
.io_out_1323(dataOut[1323]),
.io_out_1324(dataOut[1324]),
.io_out_1325(dataOut[1325]),
.io_out_1326(dataOut[1326]),
.io_out_1327(dataOut[1327]),
.io_out_1328(dataOut[1328]),
.io_out_1329(dataOut[1329]),
.io_out_1330(dataOut[1330]),
.io_out_1331(dataOut[1331]),
.io_out_1332(dataOut[1332]),
.io_out_1333(dataOut[1333]),
.io_out_1334(dataOut[1334]),
.io_out_1335(dataOut[1335]),
.io_out_1336(dataOut[1336]),
.io_out_1337(dataOut[1337]),
.io_out_1338(dataOut[1338]),
.io_out_1339(dataOut[1339]),
.io_out_1340(dataOut[1340]),
.io_out_1341(dataOut[1341]),
.io_out_1342(dataOut[1342]),
.io_out_1343(dataOut[1343]),
.io_out_1344(dataOut[1344]),
.io_out_1345(dataOut[1345]),
.io_out_1346(dataOut[1346]),
.io_out_1347(dataOut[1347]),
.io_out_1348(dataOut[1348]),
.io_out_1349(dataOut[1349]),
.io_out_1350(dataOut[1350]),
.io_out_1351(dataOut[1351]),
.io_out_1352(dataOut[1352]),
.io_out_1353(dataOut[1353]),
.io_out_1354(dataOut[1354]),
.io_out_1355(dataOut[1355]),
.io_out_1356(dataOut[1356]),
.io_out_1357(dataOut[1357]),
.io_out_1358(dataOut[1358]),
.io_out_1359(dataOut[1359]),
.io_out_1360(dataOut[1360]),
.io_out_1361(dataOut[1361]),
.io_out_1362(dataOut[1362]),
.io_out_1363(dataOut[1363]),
.io_out_1364(dataOut[1364]),
.io_out_1365(dataOut[1365]),
.io_out_1366(dataOut[1366]),
.io_out_1367(dataOut[1367]),
.io_out_1368(dataOut[1368]),
.io_out_1369(dataOut[1369]),
.io_out_1370(dataOut[1370]),
.io_out_1371(dataOut[1371]),
.io_out_1372(dataOut[1372]),
.io_out_1373(dataOut[1373]),
.io_out_1374(dataOut[1374]),
.io_out_1375(dataOut[1375]),
.io_out_1376(dataOut[1376]),
.io_out_1377(dataOut[1377]),
.io_out_1378(dataOut[1378]),
.io_out_1379(dataOut[1379]),
.io_out_1380(dataOut[1380]),
.io_out_1381(dataOut[1381]),
.io_out_1382(dataOut[1382]),
.io_out_1383(dataOut[1383]),
.io_out_1384(dataOut[1384]),
.io_out_1385(dataOut[1385]),
.io_out_1386(dataOut[1386]),
.io_out_1387(dataOut[1387]),
.io_out_1388(dataOut[1388]),
.io_out_1389(dataOut[1389]),
.io_out_1390(dataOut[1390]),
.io_out_1391(dataOut[1391]),
.io_out_1392(dataOut[1392]),
.io_out_1393(dataOut[1393]),
.io_out_1394(dataOut[1394]),
.io_out_1395(dataOut[1395]),
.io_out_1396(dataOut[1396]),
.io_out_1397(dataOut[1397]),
.io_out_1398(dataOut[1398]),
.io_out_1399(dataOut[1399]),
.io_out_1400(dataOut[1400]),
.io_out_1401(dataOut[1401]),
.io_out_1402(dataOut[1402]),
.io_out_1403(dataOut[1403]),
.io_out_1404(dataOut[1404]),
.io_out_1405(dataOut[1405]),
.io_out_1406(dataOut[1406]),
.io_out_1407(dataOut[1407]),
.io_out_1408(dataOut[1408]),
.io_out_1409(dataOut[1409]),
.io_out_1410(dataOut[1410]),
.io_out_1411(dataOut[1411]),
.io_out_1412(dataOut[1412]),
.io_out_1413(dataOut[1413]),
.io_out_1414(dataOut[1414]),
.io_out_1415(dataOut[1415]),
.io_out_1416(dataOut[1416]),
.io_out_1417(dataOut[1417]),
.io_out_1418(dataOut[1418]),
.io_out_1419(dataOut[1419]),
.io_out_1420(dataOut[1420]),
.io_out_1421(dataOut[1421]),
.io_out_1422(dataOut[1422]),
.io_out_1423(dataOut[1423]),
.io_out_1424(dataOut[1424]),
.io_out_1425(dataOut[1425]),
.io_out_1426(dataOut[1426]),
.io_out_1427(dataOut[1427]),
.io_out_1428(dataOut[1428]),
.io_out_1429(dataOut[1429]),
.io_out_1430(dataOut[1430]),
.io_out_1431(dataOut[1431]),
.io_out_1432(dataOut[1432]),
.io_out_1433(dataOut[1433]),
.io_out_1434(dataOut[1434]),
.io_out_1435(dataOut[1435]),
.io_out_1436(dataOut[1436]),
.io_out_1437(dataOut[1437]),
.io_out_1438(dataOut[1438]),
.io_out_1439(dataOut[1439]),
.io_out_1440(dataOut[1440]),
.io_out_1441(dataOut[1441]),
.io_out_1442(dataOut[1442]),
.io_out_1443(dataOut[1443]),
.io_out_1444(dataOut[1444]),
.io_out_1445(dataOut[1445]),
.io_out_1446(dataOut[1446]),
.io_out_1447(dataOut[1447]),
.io_out_1448(dataOut[1448]),
.io_out_1449(dataOut[1449]),
.io_out_1450(dataOut[1450]),
.io_out_1451(dataOut[1451]),
.io_out_1452(dataOut[1452]),
.io_out_1453(dataOut[1453]),
.io_out_1454(dataOut[1454]),
.io_out_1455(dataOut[1455]),
.io_out_1456(dataOut[1456]),
.io_out_1457(dataOut[1457]),
.io_out_1458(dataOut[1458]),
.io_out_1459(dataOut[1459]),
.io_out_1460(dataOut[1460]),
.io_out_1461(dataOut[1461]),
.io_out_1462(dataOut[1462]),
.io_out_1463(dataOut[1463]),
.io_out_1464(dataOut[1464]),
.io_out_1465(dataOut[1465]),
.io_out_1466(dataOut[1466]),
.io_out_1467(dataOut[1467]),
.io_out_1468(dataOut[1468]),
.io_out_1469(dataOut[1469]),
.io_out_1470(dataOut[1470]),
.io_out_1471(dataOut[1471]),
.io_out_1472(dataOut[1472]),
.io_out_1473(dataOut[1473]),
.io_out_1474(dataOut[1474]),
.io_out_1475(dataOut[1475]),
.io_out_1476(dataOut[1476]),
.io_out_1477(dataOut[1477]),
.io_out_1478(dataOut[1478]),
.io_out_1479(dataOut[1479]),
.io_out_1480(dataOut[1480]),
.io_out_1481(dataOut[1481]),
.io_out_1482(dataOut[1482]),
.io_out_1483(dataOut[1483]),
.io_out_1484(dataOut[1484]),
.io_out_1485(dataOut[1485]),
.io_out_1486(dataOut[1486]),
.io_out_1487(dataOut[1487]),
.io_out_1488(dataOut[1488]),
.io_out_1489(dataOut[1489]),
.io_out_1490(dataOut[1490]),
.io_out_1491(dataOut[1491]),
.io_out_1492(dataOut[1492]),
.io_out_1493(dataOut[1493]),
.io_out_1494(dataOut[1494]),
.io_out_1495(dataOut[1495]),
.io_out_1496(dataOut[1496]),
.io_out_1497(dataOut[1497]),
.io_out_1498(dataOut[1498]),
.io_out_1499(dataOut[1499]),
.io_out_1500(dataOut[1500]),
.io_out_1501(dataOut[1501]),
.io_out_1502(dataOut[1502]),
.io_out_1503(dataOut[1503]),
.io_out_1504(dataOut[1504]),
.io_out_1505(dataOut[1505]),
.io_out_1506(dataOut[1506]),
.io_out_1507(dataOut[1507]),
.io_out_1508(dataOut[1508]),
.io_out_1509(dataOut[1509]),
.io_out_1510(dataOut[1510]),
.io_out_1511(dataOut[1511]),
.io_out_1512(dataOut[1512]),
.io_out_1513(dataOut[1513]),
.io_out_1514(dataOut[1514]),
.io_out_1515(dataOut[1515]),
.io_out_1516(dataOut[1516]),
.io_out_1517(dataOut[1517]),
.io_out_1518(dataOut[1518]),
.io_out_1519(dataOut[1519]),
.io_out_1520(dataOut[1520]),
.io_out_1521(dataOut[1521]),
.io_out_1522(dataOut[1522]),
.io_out_1523(dataOut[1523]),
.io_out_1524(dataOut[1524]),
.io_out_1525(dataOut[1525]),
.io_out_1526(dataOut[1526]),
.io_out_1527(dataOut[1527]),
.io_out_1528(dataOut[1528]),
.io_out_1529(dataOut[1529]),
.io_out_1530(dataOut[1530]),
.io_out_1531(dataOut[1531]),
.io_out_1532(dataOut[1532]),
.io_out_1533(dataOut[1533]),
.io_out_1534(dataOut[1534]),
.io_out_1535(dataOut[1535]),
.io_out_1536(dataOut[1536]),
.io_out_1537(dataOut[1537]),
.io_out_1538(dataOut[1538]),
.io_out_1539(dataOut[1539]),
.io_out_1540(dataOut[1540]),
.io_out_1541(dataOut[1541]),
.io_out_1542(dataOut[1542]),
.io_out_1543(dataOut[1543]),
.io_out_1544(dataOut[1544]),
.io_out_1545(dataOut[1545]),
.io_out_1546(dataOut[1546]),
.io_out_1547(dataOut[1547]),
.io_out_1548(dataOut[1548]),
.io_out_1549(dataOut[1549]),
.io_out_1550(dataOut[1550]),
.io_out_1551(dataOut[1551]),
.io_out_1552(dataOut[1552]),
.io_out_1553(dataOut[1553]),
.io_out_1554(dataOut[1554]),
.io_out_1555(dataOut[1555]),
.io_out_1556(dataOut[1556]),
.io_out_1557(dataOut[1557]),
.io_out_1558(dataOut[1558]),
.io_out_1559(dataOut[1559]),
.io_out_1560(dataOut[1560]),
.io_out_1561(dataOut[1561]),
.io_out_1562(dataOut[1562]),
.io_out_1563(dataOut[1563]),
.io_out_1564(dataOut[1564]),
.io_out_1565(dataOut[1565]),
.io_out_1566(dataOut[1566]),
.io_out_1567(dataOut[1567]),
.io_out_1568(dataOut[1568]),
.io_out_1569(dataOut[1569]),
.io_out_1570(dataOut[1570]),
.io_out_1571(dataOut[1571]),
.io_out_1572(dataOut[1572]),
.io_out_1573(dataOut[1573]),
.io_out_1574(dataOut[1574]),
.io_out_1575(dataOut[1575]),
.io_out_1576(dataOut[1576]),
.io_out_1577(dataOut[1577]),
.io_out_1578(dataOut[1578]),
.io_out_1579(dataOut[1579]),
.io_out_1580(dataOut[1580]),
.io_out_1581(dataOut[1581]),
.io_out_1582(dataOut[1582]),
.io_out_1583(dataOut[1583]),
.io_out_1584(dataOut[1584]),
.io_out_1585(dataOut[1585]),
.io_out_1586(dataOut[1586]),
.io_out_1587(dataOut[1587]),
.io_out_1588(dataOut[1588]),
.io_out_1589(dataOut[1589]),
.io_out_1590(dataOut[1590]),
.io_out_1591(dataOut[1591]),
.io_out_1592(dataOut[1592]),
.io_out_1593(dataOut[1593]),
.io_out_1594(dataOut[1594]),
.io_out_1595(dataOut[1595]),
.io_out_1596(dataOut[1596]),
.io_out_1597(dataOut[1597]),
.io_out_1598(dataOut[1598]),
.io_out_1599(dataOut[1599]),
.io_out_1600(dataOut[1600]),
.io_out_1601(dataOut[1601]),
.io_out_1602(dataOut[1602]),
.io_out_1603(dataOut[1603]),
.io_out_1604(dataOut[1604]),
.io_out_1605(dataOut[1605]),
.io_out_1606(dataOut[1606]),
.io_out_1607(dataOut[1607]),
.io_out_1608(dataOut[1608]),
.io_out_1609(dataOut[1609]),
.io_out_1610(dataOut[1610]),
.io_out_1611(dataOut[1611]),
.io_out_1612(dataOut[1612]),
.io_out_1613(dataOut[1613]),
.io_out_1614(dataOut[1614]),
.io_out_1615(dataOut[1615]),
.io_out_1616(dataOut[1616]),
.io_out_1617(dataOut[1617]),
.io_out_1618(dataOut[1618]),
.io_out_1619(dataOut[1619]),
.io_out_1620(dataOut[1620]),
.io_out_1621(dataOut[1621]),
.io_out_1622(dataOut[1622]),
.io_out_1623(dataOut[1623]),
.io_out_1624(dataOut[1624]),
.io_out_1625(dataOut[1625]),
.io_out_1626(dataOut[1626]),
.io_out_1627(dataOut[1627]),
.io_out_1628(dataOut[1628]),
.io_out_1629(dataOut[1629]),
.io_out_1630(dataOut[1630]),
.io_out_1631(dataOut[1631]),
.io_out_1632(dataOut[1632]),
.io_out_1633(dataOut[1633]),
.io_out_1634(dataOut[1634]),
.io_out_1635(dataOut[1635]),
.io_out_1636(dataOut[1636]),
.io_out_1637(dataOut[1637]),
.io_out_1638(dataOut[1638]),
.io_out_1639(dataOut[1639]),
.io_out_1640(dataOut[1640]),
.io_out_1641(dataOut[1641]),
.io_out_1642(dataOut[1642]),
.io_out_1643(dataOut[1643]),
.io_out_1644(dataOut[1644]),
.io_out_1645(dataOut[1645]),
.io_out_1646(dataOut[1646]),
.io_out_1647(dataOut[1647]),
.io_out_1648(dataOut[1648]),
.io_out_1649(dataOut[1649]),
.io_out_1650(dataOut[1650]),
.io_out_1651(dataOut[1651]),
.io_out_1652(dataOut[1652]),
.io_out_1653(dataOut[1653]),
.io_out_1654(dataOut[1654]),
.io_out_1655(dataOut[1655]),
.io_out_1656(dataOut[1656]),
.io_out_1657(dataOut[1657]),
.io_out_1658(dataOut[1658]),
.io_out_1659(dataOut[1659]),
.io_out_1660(dataOut[1660]),
.io_out_1661(dataOut[1661]),
.io_out_1662(dataOut[1662]),
.io_out_1663(dataOut[1663]),
.io_out_1664(dataOut[1664]),
.io_out_1665(dataOut[1665]),
.io_out_1666(dataOut[1666]),
.io_out_1667(dataOut[1667]),
.io_out_1668(dataOut[1668]),
.io_out_1669(dataOut[1669]),
.io_out_1670(dataOut[1670]),
.io_out_1671(dataOut[1671]),
.io_out_1672(dataOut[1672]),
.io_out_1673(dataOut[1673]),
.io_out_1674(dataOut[1674]),
.io_out_1675(dataOut[1675]),
.io_out_1676(dataOut[1676]),
.io_out_1677(dataOut[1677]),
.io_out_1678(dataOut[1678]),
.io_out_1679(dataOut[1679]),
.io_out_1680(dataOut[1680]),
.io_out_1681(dataOut[1681]),
.io_out_1682(dataOut[1682]),
.io_out_1683(dataOut[1683]),
.io_out_1684(dataOut[1684]),
.io_out_1685(dataOut[1685]),
.io_out_1686(dataOut[1686]),
.io_out_1687(dataOut[1687]),
.io_out_1688(dataOut[1688]),
.io_out_1689(dataOut[1689]),
.io_out_1690(dataOut[1690]),
.io_out_1691(dataOut[1691]),
.io_out_1692(dataOut[1692]),
.io_out_1693(dataOut[1693]),
.io_out_1694(dataOut[1694]),
.io_out_1695(dataOut[1695]),
.io_out_1696(dataOut[1696]),
.io_out_1697(dataOut[1697]),
.io_out_1698(dataOut[1698]),
.io_out_1699(dataOut[1699]),
.io_out_1700(dataOut[1700]),
.io_out_1701(dataOut[1701]),
.io_out_1702(dataOut[1702]),
.io_out_1703(dataOut[1703]),
.io_out_1704(dataOut[1704]),
.io_out_1705(dataOut[1705]),
.io_out_1706(dataOut[1706]),
.io_out_1707(dataOut[1707]),
.io_out_1708(dataOut[1708]),
.io_out_1709(dataOut[1709]),
.io_out_1710(dataOut[1710]),
.io_out_1711(dataOut[1711]),
.io_out_1712(dataOut[1712]),
.io_out_1713(dataOut[1713]),
.io_out_1714(dataOut[1714]),
.io_out_1715(dataOut[1715]),
.io_out_1716(dataOut[1716]),
.io_out_1717(dataOut[1717]),
.io_out_1718(dataOut[1718]),
.io_out_1719(dataOut[1719]),
.io_out_1720(dataOut[1720]),
.io_out_1721(dataOut[1721]),
.io_out_1722(dataOut[1722]),
.io_out_1723(dataOut[1723]),
.io_out_1724(dataOut[1724]),
.io_out_1725(dataOut[1725]),
.io_out_1726(dataOut[1726]),
.io_out_1727(dataOut[1727]),
.io_out_1728(dataOut[1728]),
.io_out_1729(dataOut[1729]),
.io_out_1730(dataOut[1730]),
.io_out_1731(dataOut[1731]),
.io_out_1732(dataOut[1732]),
.io_out_1733(dataOut[1733]),
.io_out_1734(dataOut[1734]),
.io_out_1735(dataOut[1735]),
.io_out_1736(dataOut[1736]),
.io_out_1737(dataOut[1737]),
.io_out_1738(dataOut[1738]),
.io_out_1739(dataOut[1739]),
.io_out_1740(dataOut[1740]),
.io_out_1741(dataOut[1741]),
.io_out_1742(dataOut[1742]),
.io_out_1743(dataOut[1743]),
.io_out_1744(dataOut[1744]),
.io_out_1745(dataOut[1745]),
.io_out_1746(dataOut[1746]),
.io_out_1747(dataOut[1747]),
.io_out_1748(dataOut[1748]),
.io_out_1749(dataOut[1749]),
.io_out_1750(dataOut[1750]),
.io_out_1751(dataOut[1751]),
.io_out_1752(dataOut[1752]),
.io_out_1753(dataOut[1753]),
.io_out_1754(dataOut[1754]),
.io_out_1755(dataOut[1755]),
.io_out_1756(dataOut[1756]),
.io_out_1757(dataOut[1757]),
.io_out_1758(dataOut[1758]),
.io_out_1759(dataOut[1759]),
.io_out_1760(dataOut[1760]),
.io_out_1761(dataOut[1761]),
.io_out_1762(dataOut[1762]),
.io_out_1763(dataOut[1763]),
.io_out_1764(dataOut[1764]),
.io_out_1765(dataOut[1765]),
.io_out_1766(dataOut[1766]),
.io_out_1767(dataOut[1767]),
.io_out_1768(dataOut[1768]),
.io_out_1769(dataOut[1769]),
.io_out_1770(dataOut[1770]),
.io_out_1771(dataOut[1771]),
.io_out_1772(dataOut[1772]),
.io_out_1773(dataOut[1773]),
.io_out_1774(dataOut[1774]),
.io_out_1775(dataOut[1775]),
.io_out_1776(dataOut[1776]),
.io_out_1777(dataOut[1777]),
.io_out_1778(dataOut[1778]),
.io_out_1779(dataOut[1779]),
.io_out_1780(dataOut[1780]),
.io_out_1781(dataOut[1781]),
.io_out_1782(dataOut[1782]),
.io_out_1783(dataOut[1783]),
.io_out_1784(dataOut[1784]),
.io_out_1785(dataOut[1785]),
.io_out_1786(dataOut[1786]),
.io_out_1787(dataOut[1787]),
.io_out_1788(dataOut[1788]),
.io_out_1789(dataOut[1789]),
.io_out_1790(dataOut[1790]),
.io_out_1791(dataOut[1791]),
.io_out_1792(dataOut[1792]),
.io_out_1793(dataOut[1793]),
.io_out_1794(dataOut[1794]),
.io_out_1795(dataOut[1795]),
.io_out_1796(dataOut[1796]),
.io_out_1797(dataOut[1797]),
.io_out_1798(dataOut[1798]),
.io_out_1799(dataOut[1799]),
.io_out_1800(dataOut[1800]),
.io_out_1801(dataOut[1801]),
.io_out_1802(dataOut[1802]),
.io_out_1803(dataOut[1803]),
.io_out_1804(dataOut[1804]),
.io_out_1805(dataOut[1805]),
.io_out_1806(dataOut[1806]),
.io_out_1807(dataOut[1807]),
.io_out_1808(dataOut[1808]),
.io_out_1809(dataOut[1809]),
.io_out_1810(dataOut[1810]),
.io_out_1811(dataOut[1811]),
.io_out_1812(dataOut[1812]),
.io_out_1813(dataOut[1813]),
.io_out_1814(dataOut[1814]),
.io_out_1815(dataOut[1815]),
.io_out_1816(dataOut[1816]),
.io_out_1817(dataOut[1817]),
.io_out_1818(dataOut[1818]),
.io_out_1819(dataOut[1819]),
.io_out_1820(dataOut[1820]),
.io_out_1821(dataOut[1821]),
.io_out_1822(dataOut[1822]),
.io_out_1823(dataOut[1823]),
.io_out_1824(dataOut[1824]),
.io_out_1825(dataOut[1825]),
.io_out_1826(dataOut[1826]),
.io_out_1827(dataOut[1827]),
.io_out_1828(dataOut[1828]),
.io_out_1829(dataOut[1829]),
.io_out_1830(dataOut[1830]),
.io_out_1831(dataOut[1831]),
.io_out_1832(dataOut[1832]),
.io_out_1833(dataOut[1833]),
.io_out_1834(dataOut[1834]),
.io_out_1835(dataOut[1835]),
.io_out_1836(dataOut[1836]),
.io_out_1837(dataOut[1837]),
.io_out_1838(dataOut[1838]),
.io_out_1839(dataOut[1839]),
.io_out_1840(dataOut[1840]),
.io_out_1841(dataOut[1841]),
.io_out_1842(dataOut[1842]),
.io_out_1843(dataOut[1843]),
.io_out_1844(dataOut[1844]),
.io_out_1845(dataOut[1845]),
.io_out_1846(dataOut[1846]),
.io_out_1847(dataOut[1847]),
.io_out_1848(dataOut[1848]),
.io_out_1849(dataOut[1849]),
.io_out_1850(dataOut[1850]),
.io_out_1851(dataOut[1851]),
.io_out_1852(dataOut[1852]),
.io_out_1853(dataOut[1853]),
.io_out_1854(dataOut[1854]),
.io_out_1855(dataOut[1855]),
.io_out_1856(dataOut[1856]),
.io_out_1857(dataOut[1857]),
.io_out_1858(dataOut[1858]),
.io_out_1859(dataOut[1859]),
.io_out_1860(dataOut[1860]),
.io_out_1861(dataOut[1861]),
.io_out_1862(dataOut[1862]),
.io_out_1863(dataOut[1863]),
.io_out_1864(dataOut[1864]),
.io_out_1865(dataOut[1865]),
.io_out_1866(dataOut[1866]),
.io_out_1867(dataOut[1867]),
.io_out_1868(dataOut[1868]),
.io_out_1869(dataOut[1869]),
.io_out_1870(dataOut[1870]),
.io_out_1871(dataOut[1871]),
.io_out_1872(dataOut[1872]),
.io_out_1873(dataOut[1873]),
.io_out_1874(dataOut[1874]),
.io_out_1875(dataOut[1875]),
.io_out_1876(dataOut[1876]),
.io_out_1877(dataOut[1877]),
.io_out_1878(dataOut[1878]),
.io_out_1879(dataOut[1879]),
.io_out_1880(dataOut[1880]),
.io_out_1881(dataOut[1881]),
.io_out_1882(dataOut[1882]),
.io_out_1883(dataOut[1883]),
.io_out_1884(dataOut[1884]),
.io_out_1885(dataOut[1885]),
.io_out_1886(dataOut[1886]),
.io_out_1887(dataOut[1887]),
.io_out_1888(dataOut[1888]),
.io_out_1889(dataOut[1889]),
.io_out_1890(dataOut[1890]),
.io_out_1891(dataOut[1891]),
.io_out_1892(dataOut[1892]),
.io_out_1893(dataOut[1893]),
.io_out_1894(dataOut[1894]),
.io_out_1895(dataOut[1895]),
.io_out_1896(dataOut[1896]),
.io_out_1897(dataOut[1897]),
.io_out_1898(dataOut[1898]),
.io_out_1899(dataOut[1899]),
.io_out_1900(dataOut[1900]),
.io_out_1901(dataOut[1901]),
.io_out_1902(dataOut[1902]),
.io_out_1903(dataOut[1903]),
.io_out_1904(dataOut[1904]),
.io_out_1905(dataOut[1905]),
.io_out_1906(dataOut[1906]),
.io_out_1907(dataOut[1907]),
.io_out_1908(dataOut[1908]),
.io_out_1909(dataOut[1909]),
.io_out_1910(dataOut[1910]),
.io_out_1911(dataOut[1911]),
.io_out_1912(dataOut[1912]),
.io_out_1913(dataOut[1913]),
.io_out_1914(dataOut[1914]),
.io_out_1915(dataOut[1915]),
.io_out_1916(dataOut[1916]),
.io_out_1917(dataOut[1917]),
.io_out_1918(dataOut[1918]),
.io_out_1919(dataOut[1919]),
.io_out_1920(dataOut[1920]),
.io_out_1921(dataOut[1921]),
.io_out_1922(dataOut[1922]),
.io_out_1923(dataOut[1923]),
.io_out_1924(dataOut[1924]),
.io_out_1925(dataOut[1925]),
.io_out_1926(dataOut[1926]),
.io_out_1927(dataOut[1927]),
.io_out_1928(dataOut[1928]),
.io_out_1929(dataOut[1929]),
.io_out_1930(dataOut[1930]),
.io_out_1931(dataOut[1931]),
.io_out_1932(dataOut[1932]),
.io_out_1933(dataOut[1933]),
.io_out_1934(dataOut[1934]),
.io_out_1935(dataOut[1935]),
.io_out_1936(dataOut[1936]),
.io_out_1937(dataOut[1937]),
.io_out_1938(dataOut[1938]),
.io_out_1939(dataOut[1939]),
.io_out_1940(dataOut[1940]),
.io_out_1941(dataOut[1941]),
.io_out_1942(dataOut[1942]),
.io_out_1943(dataOut[1943]),
.io_out_1944(dataOut[1944]),
.io_out_1945(dataOut[1945]),
.io_out_1946(dataOut[1946]),
.io_out_1947(dataOut[1947]),
.io_out_1948(dataOut[1948]),
.io_out_1949(dataOut[1949]),
.io_out_1950(dataOut[1950]),
.io_out_1951(dataOut[1951]),
.io_out_1952(dataOut[1952]),
.io_out_1953(dataOut[1953]),
.io_out_1954(dataOut[1954]),
.io_out_1955(dataOut[1955]),
.io_out_1956(dataOut[1956]),
.io_out_1957(dataOut[1957]),
.io_out_1958(dataOut[1958]),
.io_out_1959(dataOut[1959]),
.io_out_1960(dataOut[1960]),
.io_out_1961(dataOut[1961]),
.io_out_1962(dataOut[1962]),
.io_out_1963(dataOut[1963]),
.io_out_1964(dataOut[1964]),
.io_out_1965(dataOut[1965]),
.io_out_1966(dataOut[1966]),
.io_out_1967(dataOut[1967]),
.io_out_1968(dataOut[1968]),
.io_out_1969(dataOut[1969]),
.io_out_1970(dataOut[1970]),
.io_out_1971(dataOut[1971]),
.io_out_1972(dataOut[1972]),
.io_out_1973(dataOut[1973]),
.io_out_1974(dataOut[1974]),
.io_out_1975(dataOut[1975]),
.io_out_1976(dataOut[1976]),
.io_out_1977(dataOut[1977]),
.io_out_1978(dataOut[1978]),
.io_out_1979(dataOut[1979]),
.io_out_1980(dataOut[1980]),
.io_out_1981(dataOut[1981]),
.io_out_1982(dataOut[1982]),
.io_out_1983(dataOut[1983]),
.io_out_1984(dataOut[1984]),
.io_out_1985(dataOut[1985]),
.io_out_1986(dataOut[1986]),
.io_out_1987(dataOut[1987]),
.io_out_1988(dataOut[1988]),
.io_out_1989(dataOut[1989]),
.io_out_1990(dataOut[1990]),
.io_out_1991(dataOut[1991]),
.io_out_1992(dataOut[1992]),
.io_out_1993(dataOut[1993]),
.io_out_1994(dataOut[1994]),
.io_out_1995(dataOut[1995]),
.io_out_1996(dataOut[1996]),
.io_out_1997(dataOut[1997]),
.io_out_1998(dataOut[1998]),
.io_out_1999(dataOut[1999]),
.io_out_2000(dataOut[2000]),
.io_out_2001(dataOut[2001]),
.io_out_2002(dataOut[2002]),
.io_out_2003(dataOut[2003]),
.io_out_2004(dataOut[2004]),
.io_out_2005(dataOut[2005]),
.io_out_2006(dataOut[2006]),
.io_out_2007(dataOut[2007]),
.io_out_2008(dataOut[2008]),
.io_out_2009(dataOut[2009]),
.io_out_2010(dataOut[2010]),
.io_out_2011(dataOut[2011]),
.io_out_2012(dataOut[2012]),
.io_out_2013(dataOut[2013]),
.io_out_2014(dataOut[2014]),
.io_out_2015(dataOut[2015]),
.io_out_2016(dataOut[2016]),
.io_out_2017(dataOut[2017]),
.io_out_2018(dataOut[2018]),
.io_out_2019(dataOut[2019]),
.io_out_2020(dataOut[2020]),
.io_out_2021(dataOut[2021]),
.io_out_2022(dataOut[2022]),
.io_out_2023(dataOut[2023]),
.io_out_2024(dataOut[2024]),
.io_out_2025(dataOut[2025]),
.io_out_2026(dataOut[2026]),
.io_out_2027(dataOut[2027]),
.io_out_2028(dataOut[2028]),
.io_out_2029(dataOut[2029]),
.io_out_2030(dataOut[2030]),
.io_out_2031(dataOut[2031]),
.io_out_2032(dataOut[2032]),
.io_out_2033(dataOut[2033]),
.io_out_2034(dataOut[2034]),
.io_out_2035(dataOut[2035]),
.io_out_2036(dataOut[2036]),
.io_out_2037(dataOut[2037]),
.io_out_2038(dataOut[2038]),
.io_out_2039(dataOut[2039]),
.io_out_2040(dataOut[2040]),
.io_out_2041(dataOut[2041]),
.io_out_2042(dataOut[2042]),
.io_out_2043(dataOut[2043]),
.io_out_2044(dataOut[2044]),
.io_out_2045(dataOut[2045]),
.io_out_2046(dataOut[2046]),
.io_out_2047(dataOut[2047]),
.io_out_2048(dataOut[2048]),
.io_out_2049(dataOut[2049]),
.io_out_2050(dataOut[2050]),
.io_out_2051(dataOut[2051]),
.io_out_2052(dataOut[2052]),
.io_out_2053(dataOut[2053]),
.io_out_2054(dataOut[2054]),
.io_out_2055(dataOut[2055]),
.io_out_2056(dataOut[2056]),
.io_out_2057(dataOut[2057]),
.io_out_2058(dataOut[2058]),
.io_out_2059(dataOut[2059]),
.io_out_2060(dataOut[2060]),
.io_out_2061(dataOut[2061]),
.io_out_2062(dataOut[2062]),
.io_out_2063(dataOut[2063]),
.io_out_2064(dataOut[2064]),
.io_out_2065(dataOut[2065]),
.io_out_2066(dataOut[2066]),
.io_out_2067(dataOut[2067]),
.io_out_2068(dataOut[2068]),
.io_out_2069(dataOut[2069]),
.io_out_2070(dataOut[2070]),
.io_out_2071(dataOut[2071]),
.io_out_2072(dataOut[2072]),
.io_out_2073(dataOut[2073]),
.io_out_2074(dataOut[2074]),
.io_out_2075(dataOut[2075]),
.io_out_2076(dataOut[2076]),
.io_out_2077(dataOut[2077]),
.io_out_2078(dataOut[2078]),
.io_out_2079(dataOut[2079]),
.io_out_2080(dataOut[2080]),
.io_out_2081(dataOut[2081]),
.io_out_2082(dataOut[2082]),
.io_out_2083(dataOut[2083]),
.io_out_2084(dataOut[2084]),
.io_out_2085(dataOut[2085]),
.io_out_2086(dataOut[2086]),
.io_out_2087(dataOut[2087]),
.io_out_2088(dataOut[2088]),
.io_out_2089(dataOut[2089]),
.io_out_2090(dataOut[2090]),
.io_out_2091(dataOut[2091]),
.io_out_2092(dataOut[2092]),
.io_out_2093(dataOut[2093]),
.io_out_2094(dataOut[2094]),
.io_out_2095(dataOut[2095]),
.io_out_2096(dataOut[2096]),
.io_out_2097(dataOut[2097]),
.io_out_2098(dataOut[2098]),
.io_out_2099(dataOut[2099]),
.io_out_2100(dataOut[2100]),
.io_out_2101(dataOut[2101]),
.io_out_2102(dataOut[2102]),
.io_out_2103(dataOut[2103]),
.io_out_2104(dataOut[2104]),
.io_out_2105(dataOut[2105]),
.io_out_2106(dataOut[2106]),
.io_out_2107(dataOut[2107]),
.io_out_2108(dataOut[2108]),
.io_out_2109(dataOut[2109]),
.io_out_2110(dataOut[2110]),
.io_out_2111(dataOut[2111]),
.io_out_2112(dataOut[2112]),
.io_out_2113(dataOut[2113]),
.io_out_2114(dataOut[2114]),
.io_out_2115(dataOut[2115]),
.io_out_2116(dataOut[2116]),
.io_out_2117(dataOut[2117]),
.io_out_2118(dataOut[2118]),
.io_out_2119(dataOut[2119]),
.io_out_2120(dataOut[2120]),
.io_out_2121(dataOut[2121]),
.io_out_2122(dataOut[2122]),
.io_out_2123(dataOut[2123]),
.io_out_2124(dataOut[2124]),
.io_out_2125(dataOut[2125]),
.io_out_2126(dataOut[2126]),
.io_out_2127(dataOut[2127]),
.io_out_2128(dataOut[2128]),
.io_out_2129(dataOut[2129]),
.io_out_2130(dataOut[2130]),
.io_out_2131(dataOut[2131]),
.io_out_2132(dataOut[2132]),
.io_out_2133(dataOut[2133]),
.io_out_2134(dataOut[2134]),
.io_out_2135(dataOut[2135]),
.io_out_2136(dataOut[2136]),
.io_out_2137(dataOut[2137]),
.io_out_2138(dataOut[2138]),
.io_out_2139(dataOut[2139]),
.io_out_2140(dataOut[2140]),
.io_out_2141(dataOut[2141]),
.io_out_2142(dataOut[2142]),
.io_out_2143(dataOut[2143]),
.io_out_2144(dataOut[2144]),
.io_out_2145(dataOut[2145]),
.io_out_2146(dataOut[2146]),
.io_out_2147(dataOut[2147]),
.io_out_2148(dataOut[2148]),
.io_out_2149(dataOut[2149]),
.io_out_2150(dataOut[2150]),
.io_out_2151(dataOut[2151]),
.io_out_2152(dataOut[2152]),
.io_out_2153(dataOut[2153]),
.io_out_2154(dataOut[2154]),
.io_out_2155(dataOut[2155]),
.io_out_2156(dataOut[2156]),
.io_out_2157(dataOut[2157]),
.io_out_2158(dataOut[2158]),
.io_out_2159(dataOut[2159]),
.io_out_2160(dataOut[2160]),
.io_out_2161(dataOut[2161]),
.io_out_2162(dataOut[2162]),
.io_out_2163(dataOut[2163]),
.io_out_2164(dataOut[2164]),
.io_out_2165(dataOut[2165]),
.io_out_2166(dataOut[2166]),
.io_out_2167(dataOut[2167]),
.io_out_2168(dataOut[2168]),
.io_out_2169(dataOut[2169]),
.io_out_2170(dataOut[2170]),
.io_out_2171(dataOut[2171]),
.io_out_2172(dataOut[2172]),
.io_out_2173(dataOut[2173]),
.io_out_2174(dataOut[2174]),
.io_out_2175(dataOut[2175]),
.io_out_2176(dataOut[2176]),
.io_out_2177(dataOut[2177]),
.io_out_2178(dataOut[2178]),
.io_out_2179(dataOut[2179]),
.io_out_2180(dataOut[2180]),
.io_out_2181(dataOut[2181]),
.io_out_2182(dataOut[2182]),
.io_out_2183(dataOut[2183]),
.io_out_2184(dataOut[2184]),
.io_out_2185(dataOut[2185]),
.io_out_2186(dataOut[2186]),
.io_out_2187(dataOut[2187]),
.io_out_2188(dataOut[2188]),
.io_out_2189(dataOut[2189]),
.io_out_2190(dataOut[2190]),
.io_out_2191(dataOut[2191]),
.io_out_2192(dataOut[2192]),
.io_out_2193(dataOut[2193]),
.io_out_2194(dataOut[2194]),
.io_out_2195(dataOut[2195]),
.io_out_2196(dataOut[2196]),
.io_out_2197(dataOut[2197]),
.io_out_2198(dataOut[2198]),
.io_out_2199(dataOut[2199]),
.io_out_2200(dataOut[2200]),
.io_out_2201(dataOut[2201]),
.io_out_2202(dataOut[2202]),
.io_out_2203(dataOut[2203]),
.io_out_2204(dataOut[2204]),
.io_out_2205(dataOut[2205]),
.io_out_2206(dataOut[2206]),
.io_out_2207(dataOut[2207]),
.io_out_2208(dataOut[2208]),
.io_out_2209(dataOut[2209]),
.io_out_2210(dataOut[2210]),
.io_out_2211(dataOut[2211]),
.io_out_2212(dataOut[2212]),
.io_out_2213(dataOut[2213]),
.io_out_2214(dataOut[2214]),
.io_out_2215(dataOut[2215]),
.io_out_2216(dataOut[2216]),
.io_out_2217(dataOut[2217]),
.io_out_2218(dataOut[2218]),
.io_out_2219(dataOut[2219]),
.io_out_2220(dataOut[2220]),
.io_out_2221(dataOut[2221]),
.io_out_2222(dataOut[2222]),
.io_out_2223(dataOut[2223]),
.io_out_2224(dataOut[2224]),
.io_out_2225(dataOut[2225]),
.io_out_2226(dataOut[2226]),
.io_out_2227(dataOut[2227]),
.io_out_2228(dataOut[2228]),
.io_out_2229(dataOut[2229]),
.io_out_2230(dataOut[2230]),
.io_out_2231(dataOut[2231]),
.io_out_2232(dataOut[2232]),
.io_out_2233(dataOut[2233]),
.io_out_2234(dataOut[2234]),
.io_out_2235(dataOut[2235]),
.io_out_2236(dataOut[2236]),
.io_out_2237(dataOut[2237]),
.io_out_2238(dataOut[2238]),
.io_out_2239(dataOut[2239]),
.io_out_2240(dataOut[2240]),
.io_out_2241(dataOut[2241]),
.io_out_2242(dataOut[2242]),
.io_out_2243(dataOut[2243]),
.io_out_2244(dataOut[2244]),
.io_out_2245(dataOut[2245]),
.io_out_2246(dataOut[2246]),
.io_out_2247(dataOut[2247]),
.io_out_2248(dataOut[2248]),
.io_out_2249(dataOut[2249]),
.io_out_2250(dataOut[2250]),
.io_out_2251(dataOut[2251]),
.io_out_2252(dataOut[2252]),
.io_out_2253(dataOut[2253]),
.io_out_2254(dataOut[2254]),
.io_out_2255(dataOut[2255]),
.io_out_2256(dataOut[2256]),
.io_out_2257(dataOut[2257]),
.io_out_2258(dataOut[2258]),
.io_out_2259(dataOut[2259]),
.io_out_2260(dataOut[2260]),
.io_out_2261(dataOut[2261]),
.io_out_2262(dataOut[2262]),
.io_out_2263(dataOut[2263]),
.io_out_2264(dataOut[2264]),
.io_out_2265(dataOut[2265]),
.io_out_2266(dataOut[2266]),
.io_out_2267(dataOut[2267]),
.io_out_2268(dataOut[2268]),
.io_out_2269(dataOut[2269]),
.io_out_2270(dataOut[2270]),
.io_out_2271(dataOut[2271]),
.io_out_2272(dataOut[2272]),
.io_out_2273(dataOut[2273]),
.io_out_2274(dataOut[2274]),
.io_out_2275(dataOut[2275]),
.io_out_2276(dataOut[2276]),
.io_out_2277(dataOut[2277]),
.io_out_2278(dataOut[2278]),
.io_out_2279(dataOut[2279]),
.io_out_2280(dataOut[2280]),
.io_out_2281(dataOut[2281]),
.io_out_2282(dataOut[2282]),
.io_out_2283(dataOut[2283]),
.io_out_2284(dataOut[2284]),
.io_out_2285(dataOut[2285]),
.io_out_2286(dataOut[2286]),
.io_out_2287(dataOut[2287]),
.io_out_2288(dataOut[2288]),
.io_out_2289(dataOut[2289]),
.io_out_2290(dataOut[2290]),
.io_out_2291(dataOut[2291]),
.io_out_2292(dataOut[2292]),
.io_out_2293(dataOut[2293]),
.io_out_2294(dataOut[2294]),
.io_out_2295(dataOut[2295]),
.io_out_2296(dataOut[2296]),
.io_out_2297(dataOut[2297]),
.io_out_2298(dataOut[2298]),
.io_out_2299(dataOut[2299]),
.io_out_2300(dataOut[2300]),
.io_out_2301(dataOut[2301]),
.io_out_2302(dataOut[2302]),
.io_out_2303(dataOut[2303]),
.io_out_2304(dataOut[2304]),
.io_out_2305(dataOut[2305]),
.io_out_2306(dataOut[2306]),
.io_out_2307(dataOut[2307]),
.io_out_2308(dataOut[2308]),
.io_out_2309(dataOut[2309]),
.io_out_2310(dataOut[2310]),
.io_out_2311(dataOut[2311]),
.io_out_2312(dataOut[2312]),
.io_out_2313(dataOut[2313]),
.io_out_2314(dataOut[2314]),
.io_out_2315(dataOut[2315]),
.io_out_2316(dataOut[2316]),
.io_out_2317(dataOut[2317]),
.io_out_2318(dataOut[2318]),
.io_out_2319(dataOut[2319]),
.io_out_2320(dataOut[2320]),
.io_out_2321(dataOut[2321]),
.io_out_2322(dataOut[2322]),
.io_out_2323(dataOut[2323]),
.io_out_2324(dataOut[2324]),
.io_out_2325(dataOut[2325]),
.io_out_2326(dataOut[2326]),
.io_out_2327(dataOut[2327]),
.io_out_2328(dataOut[2328]),
.io_out_2329(dataOut[2329]),
.io_out_2330(dataOut[2330]),
.io_out_2331(dataOut[2331]),
.io_out_2332(dataOut[2332]),
.io_out_2333(dataOut[2333]),
.io_out_2334(dataOut[2334]),
.io_out_2335(dataOut[2335]),
.io_out_2336(dataOut[2336]),
.io_out_2337(dataOut[2337]),
.io_out_2338(dataOut[2338]),
.io_out_2339(dataOut[2339]),
.io_out_2340(dataOut[2340]),
.io_out_2341(dataOut[2341]),
.io_out_2342(dataOut[2342]),
.io_out_2343(dataOut[2343]),
.io_out_2344(dataOut[2344]),
.io_out_2345(dataOut[2345]),
.io_out_2346(dataOut[2346]),
.io_out_2347(dataOut[2347]),
.io_out_2348(dataOut[2348]),
.io_out_2349(dataOut[2349]),
.io_out_2350(dataOut[2350]),
.io_out_2351(dataOut[2351]),
.io_out_2352(dataOut[2352]),
.io_out_2353(dataOut[2353]),
.io_out_2354(dataOut[2354]),
.io_out_2355(dataOut[2355]),
.io_out_2356(dataOut[2356]),
.io_out_2357(dataOut[2357]),
.io_out_2358(dataOut[2358]),
.io_out_2359(dataOut[2359]),
.io_out_2360(dataOut[2360]),
.io_out_2361(dataOut[2361]),
.io_out_2362(dataOut[2362]),
.io_out_2363(dataOut[2363]),
.io_out_2364(dataOut[2364]),
.io_out_2365(dataOut[2365]),
.io_out_2366(dataOut[2366]),
.io_out_2367(dataOut[2367]),
.io_out_2368(dataOut[2368]),
.io_out_2369(dataOut[2369]),
.io_out_2370(dataOut[2370]),
.io_out_2371(dataOut[2371]),
.io_out_2372(dataOut[2372]),
.io_out_2373(dataOut[2373]),
.io_out_2374(dataOut[2374]),
.io_out_2375(dataOut[2375]),
.io_out_2376(dataOut[2376]),
.io_out_2377(dataOut[2377]),
.io_out_2378(dataOut[2378]),
.io_out_2379(dataOut[2379]),
.io_out_2380(dataOut[2380]),
.io_out_2381(dataOut[2381]),
.io_out_2382(dataOut[2382]),
.io_out_2383(dataOut[2383]),
.io_out_2384(dataOut[2384]),
.io_out_2385(dataOut[2385]),
.io_out_2386(dataOut[2386]),
.io_out_2387(dataOut[2387]),
.io_out_2388(dataOut[2388]),
.io_out_2389(dataOut[2389]),
.io_out_2390(dataOut[2390]),
.io_out_2391(dataOut[2391]),
.io_out_2392(dataOut[2392]),
.io_out_2393(dataOut[2393]),
.io_out_2394(dataOut[2394]),
.io_out_2395(dataOut[2395]),
.io_out_2396(dataOut[2396]),
.io_out_2397(dataOut[2397]),
.io_out_2398(dataOut[2398]),
.io_out_2399(dataOut[2399]),
.io_out_2400(dataOut[2400]),
.io_out_2401(dataOut[2401]),
.io_out_2402(dataOut[2402]),
.io_out_2403(dataOut[2403]),
.io_out_2404(dataOut[2404]),
.io_out_2405(dataOut[2405]),
.io_out_2406(dataOut[2406]),
.io_out_2407(dataOut[2407]),
.io_out_2408(dataOut[2408]),
.io_out_2409(dataOut[2409]),
.io_out_2410(dataOut[2410]),
.io_out_2411(dataOut[2411]),
.io_out_2412(dataOut[2412]),
.io_out_2413(dataOut[2413]),
.io_out_2414(dataOut[2414]),
.io_out_2415(dataOut[2415]),
.io_out_2416(dataOut[2416]),
.io_out_2417(dataOut[2417]),
.io_out_2418(dataOut[2418]),
.io_out_2419(dataOut[2419]),
.io_out_2420(dataOut[2420]),
.io_out_2421(dataOut[2421]),
.io_out_2422(dataOut[2422]),
.io_out_2423(dataOut[2423]),
.io_out_2424(dataOut[2424]),
.io_out_2425(dataOut[2425]),
.io_out_2426(dataOut[2426]),
.io_out_2427(dataOut[2427]),
.io_out_2428(dataOut[2428]),
.io_out_2429(dataOut[2429]),
.io_out_2430(dataOut[2430]),
.io_out_2431(dataOut[2431]),
.io_out_2432(dataOut[2432]),
.io_out_2433(dataOut[2433]),
.io_out_2434(dataOut[2434]),
.io_out_2435(dataOut[2435]),
.io_out_2436(dataOut[2436]),
.io_out_2437(dataOut[2437]),
.io_out_2438(dataOut[2438]),
.io_out_2439(dataOut[2439]),
.io_out_2440(dataOut[2440]),
.io_out_2441(dataOut[2441]),
.io_out_2442(dataOut[2442]),
.io_out_2443(dataOut[2443]),
.io_out_2444(dataOut[2444]),
.io_out_2445(dataOut[2445]),
.io_out_2446(dataOut[2446]),
.io_out_2447(dataOut[2447]),
.io_out_2448(dataOut[2448]),
.io_out_2449(dataOut[2449]),
.io_out_2450(dataOut[2450]),
.io_out_2451(dataOut[2451]),
.io_out_2452(dataOut[2452]),
.io_out_2453(dataOut[2453]),
.io_out_2454(dataOut[2454]),
.io_out_2455(dataOut[2455]),
.io_out_2456(dataOut[2456]),
.io_out_2457(dataOut[2457]),
.io_out_2458(dataOut[2458]),
.io_out_2459(dataOut[2459]),
.io_out_2460(dataOut[2460]),
.io_out_2461(dataOut[2461]),
.io_out_2462(dataOut[2462]),
.io_out_2463(dataOut[2463]),
.io_out_2464(dataOut[2464]),
.io_out_2465(dataOut[2465]),
.io_out_2466(dataOut[2466]),
.io_out_2467(dataOut[2467]),
.io_out_2468(dataOut[2468]),
.io_out_2469(dataOut[2469]),
.io_out_2470(dataOut[2470]),
.io_out_2471(dataOut[2471]),
.io_out_2472(dataOut[2472]),
.io_out_2473(dataOut[2473]),
.io_out_2474(dataOut[2474]),
.io_out_2475(dataOut[2475]),
.io_out_2476(dataOut[2476]),
.io_out_2477(dataOut[2477]),
.io_out_2478(dataOut[2478]),
.io_out_2479(dataOut[2479]),
.io_out_2480(dataOut[2480]),
.io_out_2481(dataOut[2481]),
.io_out_2482(dataOut[2482]),
.io_out_2483(dataOut[2483]),
.io_out_2484(dataOut[2484]),
.io_out_2485(dataOut[2485]),
.io_out_2486(dataOut[2486]),
.io_out_2487(dataOut[2487]),
.io_out_2488(dataOut[2488]),
.io_out_2489(dataOut[2489]),
.io_out_2490(dataOut[2490]),
.io_out_2491(dataOut[2491]),
.io_out_2492(dataOut[2492]),
.io_out_2493(dataOut[2493]),
.io_out_2494(dataOut[2494]),
.io_out_2495(dataOut[2495]),
.io_out_2496(dataOut[2496]),
.io_out_2497(dataOut[2497]),
.io_out_2498(dataOut[2498]),
.io_out_2499(dataOut[2499]),
.io_out_2500(dataOut[2500]),
.io_out_2501(dataOut[2501]),
.io_out_2502(dataOut[2502]),
.io_out_2503(dataOut[2503]),
.io_out_2504(dataOut[2504]),
.io_out_2505(dataOut[2505]),
.io_out_2506(dataOut[2506]),
.io_out_2507(dataOut[2507]),
.io_out_2508(dataOut[2508]),
.io_out_2509(dataOut[2509]),
.io_out_2510(dataOut[2510]),
.io_out_2511(dataOut[2511]),
.io_out_2512(dataOut[2512]),
.io_out_2513(dataOut[2513]),
.io_out_2514(dataOut[2514]),
.io_out_2515(dataOut[2515]),
.io_out_2516(dataOut[2516]),
.io_out_2517(dataOut[2517]),
.io_out_2518(dataOut[2518]),
.io_out_2519(dataOut[2519]),
.io_out_2520(dataOut[2520]),
.io_out_2521(dataOut[2521]),
.io_out_2522(dataOut[2522]),
.io_out_2523(dataOut[2523]),
.io_out_2524(dataOut[2524]),
.io_out_2525(dataOut[2525]),
.io_out_2526(dataOut[2526]),
.io_out_2527(dataOut[2527]),
.io_out_2528(dataOut[2528]),
.io_out_2529(dataOut[2529]),
.io_out_2530(dataOut[2530]),
.io_out_2531(dataOut[2531]),
.io_out_2532(dataOut[2532]),
.io_out_2533(dataOut[2533]),
.io_out_2534(dataOut[2534]),
.io_out_2535(dataOut[2535]),
.io_out_2536(dataOut[2536]),
.io_out_2537(dataOut[2537]),
.io_out_2538(dataOut[2538]),
.io_out_2539(dataOut[2539]),
.io_out_2540(dataOut[2540]),
.io_out_2541(dataOut[2541]),
.io_out_2542(dataOut[2542]),
.io_out_2543(dataOut[2543]),
.io_out_2544(dataOut[2544]),
.io_out_2545(dataOut[2545]),
.io_out_2546(dataOut[2546]),
.io_out_2547(dataOut[2547]),
.io_out_2548(dataOut[2548]),
.io_out_2549(dataOut[2549]),
.io_out_2550(dataOut[2550]),
.io_out_2551(dataOut[2551]),
.io_out_2552(dataOut[2552]),
.io_out_2553(dataOut[2553]),
.io_out_2554(dataOut[2554]),
.io_out_2555(dataOut[2555]),
.io_out_2556(dataOut[2556]),
.io_out_2557(dataOut[2557]),
.io_out_2558(dataOut[2558]),
.io_out_2559(dataOut[2559]),
.io_out_2560(dataOut[2560]),
.io_out_2561(dataOut[2561]),
.io_out_2562(dataOut[2562]),
.io_out_2563(dataOut[2563]),
.io_out_2564(dataOut[2564]),
.io_out_2565(dataOut[2565]),
.io_out_2566(dataOut[2566]),
.io_out_2567(dataOut[2567]),
.io_out_2568(dataOut[2568]),
.io_out_2569(dataOut[2569]),
.io_out_2570(dataOut[2570]),
.io_out_2571(dataOut[2571]),
.io_out_2572(dataOut[2572]),
.io_out_2573(dataOut[2573]),
.io_out_2574(dataOut[2574]),
.io_out_2575(dataOut[2575]),
.io_out_2576(dataOut[2576]),
.io_out_2577(dataOut[2577]),
.io_out_2578(dataOut[2578]),
.io_out_2579(dataOut[2579]),
.io_out_2580(dataOut[2580]),
.io_out_2581(dataOut[2581]),
.io_out_2582(dataOut[2582]),
.io_out_2583(dataOut[2583]),
.io_out_2584(dataOut[2584]),
.io_out_2585(dataOut[2585]),
.io_out_2586(dataOut[2586]),
.io_out_2587(dataOut[2587]),
.io_out_2588(dataOut[2588]),
.io_out_2589(dataOut[2589]),
.io_out_2590(dataOut[2590]),
.io_out_2591(dataOut[2591]),
.io_out_2592(dataOut[2592]),
.io_out_2593(dataOut[2593]),
.io_out_2594(dataOut[2594]),
.io_out_2595(dataOut[2595]),
.io_out_2596(dataOut[2596]),
.io_out_2597(dataOut[2597]),
.io_out_2598(dataOut[2598]),
.io_out_2599(dataOut[2599]),
.io_out_2600(dataOut[2600]),
.io_out_2601(dataOut[2601]),
.io_out_2602(dataOut[2602]),
.io_out_2603(dataOut[2603]),
.io_out_2604(dataOut[2604]),
.io_out_2605(dataOut[2605]),
.io_out_2606(dataOut[2606]),
.io_out_2607(dataOut[2607]),
.io_out_2608(dataOut[2608]),
.io_out_2609(dataOut[2609]),
.io_out_2610(dataOut[2610]),
.io_out_2611(dataOut[2611]),
.io_out_2612(dataOut[2612]),
.io_out_2613(dataOut[2613]),
.io_out_2614(dataOut[2614]),
.io_out_2615(dataOut[2615]),
.io_out_2616(dataOut[2616]),
.io_out_2617(dataOut[2617]),
.io_out_2618(dataOut[2618]),
.io_out_2619(dataOut[2619]),
.io_out_2620(dataOut[2620]),
.io_out_2621(dataOut[2621]),
.io_out_2622(dataOut[2622]),
.io_out_2623(dataOut[2623]),
.io_out_2624(dataOut[2624]),
.io_out_2625(dataOut[2625]),
.io_out_2626(dataOut[2626]),
.io_out_2627(dataOut[2627]),
.io_out_2628(dataOut[2628]),
.io_out_2629(dataOut[2629]),
.io_out_2630(dataOut[2630]),
.io_out_2631(dataOut[2631]),
.io_out_2632(dataOut[2632]),
.io_out_2633(dataOut[2633]),
.io_out_2634(dataOut[2634]),
.io_out_2635(dataOut[2635]),
.io_out_2636(dataOut[2636]),
.io_out_2637(dataOut[2637]),
.io_out_2638(dataOut[2638]),
.io_out_2639(dataOut[2639]),
.io_out_2640(dataOut[2640]),
.io_out_2641(dataOut[2641]),
.io_out_2642(dataOut[2642]),
.io_out_2643(dataOut[2643]),
.io_out_2644(dataOut[2644]),
.io_out_2645(dataOut[2645]),
.io_out_2646(dataOut[2646]),
.io_out_2647(dataOut[2647]),
.io_out_2648(dataOut[2648]),
.io_out_2649(dataOut[2649]),
.io_out_2650(dataOut[2650]),
.io_out_2651(dataOut[2651]),
.io_out_2652(dataOut[2652]),
.io_out_2653(dataOut[2653]),
.io_out_2654(dataOut[2654]),
.io_out_2655(dataOut[2655]),
.io_out_2656(dataOut[2656]),
.io_out_2657(dataOut[2657]),
.io_out_2658(dataOut[2658]),
.io_out_2659(dataOut[2659]),
.io_out_2660(dataOut[2660]),
.io_out_2661(dataOut[2661]),
.io_out_2662(dataOut[2662]),
.io_out_2663(dataOut[2663]),
.io_out_2664(dataOut[2664]),
.io_out_2665(dataOut[2665]),
.io_out_2666(dataOut[2666]),
.io_out_2667(dataOut[2667]),
.io_out_2668(dataOut[2668]),
.io_out_2669(dataOut[2669]),
.io_out_2670(dataOut[2670]),
.io_out_2671(dataOut[2671]),
.io_out_2672(dataOut[2672]),
.io_out_2673(dataOut[2673]),
.io_out_2674(dataOut[2674]),
.io_out_2675(dataOut[2675]),
.io_out_2676(dataOut[2676]),
.io_out_2677(dataOut[2677]),
.io_out_2678(dataOut[2678]),
.io_out_2679(dataOut[2679]),
.io_out_2680(dataOut[2680]),
.io_out_2681(dataOut[2681]),
.io_out_2682(dataOut[2682]),
.io_out_2683(dataOut[2683]),
.io_out_2684(dataOut[2684]),
.io_out_2685(dataOut[2685]),
.io_out_2686(dataOut[2686]),
.io_out_2687(dataOut[2687]),
.io_out_2688(dataOut[2688]),
.io_out_2689(dataOut[2689]),
.io_out_2690(dataOut[2690]),
.io_out_2691(dataOut[2691]),
.io_out_2692(dataOut[2692]),
.io_out_2693(dataOut[2693]),
.io_out_2694(dataOut[2694]),
.io_out_2695(dataOut[2695]),
.io_out_2696(dataOut[2696]),
.io_out_2697(dataOut[2697]),
.io_out_2698(dataOut[2698]),
.io_out_2699(dataOut[2699]),
.io_out_2700(dataOut[2700]),
.io_out_2701(dataOut[2701]),
.io_out_2702(dataOut[2702]),
.io_out_2703(dataOut[2703]),
.io_out_2704(dataOut[2704]),
.io_out_2705(dataOut[2705]),
.io_out_2706(dataOut[2706]),
.io_out_2707(dataOut[2707]),
.io_out_2708(dataOut[2708]),
.io_out_2709(dataOut[2709]),
.io_out_2710(dataOut[2710]),
.io_out_2711(dataOut[2711]),
.io_out_2712(dataOut[2712]),
.io_out_2713(dataOut[2713]),
.io_out_2714(dataOut[2714]),
.io_out_2715(dataOut[2715]),
.io_out_2716(dataOut[2716]),
.io_out_2717(dataOut[2717]),
.io_out_2718(dataOut[2718]),
.io_out_2719(dataOut[2719]),
.io_out_2720(dataOut[2720]),
.io_out_2721(dataOut[2721]),
.io_out_2722(dataOut[2722]),
.io_out_2723(dataOut[2723]),
.io_out_2724(dataOut[2724]),
.io_out_2725(dataOut[2725]),
.io_out_2726(dataOut[2726]),
.io_out_2727(dataOut[2727]),
.io_out_2728(dataOut[2728]),
.io_out_2729(dataOut[2729]),
.io_out_2730(dataOut[2730]),
.io_out_2731(dataOut[2731]),
.io_out_2732(dataOut[2732]),
.io_out_2733(dataOut[2733]),
.io_out_2734(dataOut[2734]),
.io_out_2735(dataOut[2735]),
.io_out_2736(dataOut[2736]),
.io_out_2737(dataOut[2737]),
.io_out_2738(dataOut[2738]),
.io_out_2739(dataOut[2739]),
.io_out_2740(dataOut[2740]),
.io_out_2741(dataOut[2741]),
.io_out_2742(dataOut[2742]),
.io_out_2743(dataOut[2743]),
.io_out_2744(dataOut[2744]),
.io_out_2745(dataOut[2745]),
.io_out_2746(dataOut[2746]),
.io_out_2747(dataOut[2747]),
.io_out_2748(dataOut[2748]),
.io_out_2749(dataOut[2749]),
.io_out_2750(dataOut[2750]),
.io_out_2751(dataOut[2751]),
.io_out_2752(dataOut[2752]),
.io_out_2753(dataOut[2753]),
.io_out_2754(dataOut[2754]),
.io_out_2755(dataOut[2755]),
.io_out_2756(dataOut[2756]),
.io_out_2757(dataOut[2757]),
.io_out_2758(dataOut[2758]),
.io_out_2759(dataOut[2759]),
.io_out_2760(dataOut[2760]),
.io_out_2761(dataOut[2761]),
.io_out_2762(dataOut[2762]),
.io_out_2763(dataOut[2763]),
.io_out_2764(dataOut[2764]),
.io_out_2765(dataOut[2765]),
.io_out_2766(dataOut[2766]),
.io_out_2767(dataOut[2767]),
.io_out_2768(dataOut[2768]),
.io_out_2769(dataOut[2769]),
.io_out_2770(dataOut[2770]),
.io_out_2771(dataOut[2771]),
.io_out_2772(dataOut[2772]),
.io_out_2773(dataOut[2773]),
.io_out_2774(dataOut[2774]),
.io_out_2775(dataOut[2775]),
.io_out_2776(dataOut[2776]),
.io_out_2777(dataOut[2777]),
.io_out_2778(dataOut[2778]),
.io_out_2779(dataOut[2779]),
.io_out_2780(dataOut[2780]),
.io_out_2781(dataOut[2781]),
.io_out_2782(dataOut[2782]),
.io_out_2783(dataOut[2783]),
.io_out_2784(dataOut[2784]),
.io_out_2785(dataOut[2785]),
.io_out_2786(dataOut[2786]),
.io_out_2787(dataOut[2787]),
.io_out_2788(dataOut[2788]),
.io_out_2789(dataOut[2789]),
.io_out_2790(dataOut[2790]),
.io_out_2791(dataOut[2791]),
.io_out_2792(dataOut[2792]),
.io_out_2793(dataOut[2793]),
.io_out_2794(dataOut[2794]),
.io_out_2795(dataOut[2795]),
.io_out_2796(dataOut[2796]),
.io_out_2797(dataOut[2797]),
.io_out_2798(dataOut[2798]),
.io_out_2799(dataOut[2799]),
.io_out_2800(dataOut[2800]),
.io_out_2801(dataOut[2801]),
.io_out_2802(dataOut[2802]),
.io_out_2803(dataOut[2803]),
.io_out_2804(dataOut[2804]),
.io_out_2805(dataOut[2805]),
.io_out_2806(dataOut[2806]),
.io_out_2807(dataOut[2807]),
.io_out_2808(dataOut[2808]),
.io_out_2809(dataOut[2809]),
.io_out_2810(dataOut[2810]),
.io_out_2811(dataOut[2811]),
.io_out_2812(dataOut[2812]),
.io_out_2813(dataOut[2813]),
.io_out_2814(dataOut[2814]),
.io_out_2815(dataOut[2815]),
.io_out_2816(dataOut[2816]),
.io_out_2817(dataOut[2817]),
.io_out_2818(dataOut[2818]),
.io_out_2819(dataOut[2819]),
.io_out_2820(dataOut[2820]),
.io_out_2821(dataOut[2821]),
.io_out_2822(dataOut[2822]),
.io_out_2823(dataOut[2823]),
.io_out_2824(dataOut[2824]),
.io_out_2825(dataOut[2825]),
.io_out_2826(dataOut[2826]),
.io_out_2827(dataOut[2827]),
.io_out_2828(dataOut[2828]),
.io_out_2829(dataOut[2829]),
.io_out_2830(dataOut[2830]),
.io_out_2831(dataOut[2831]),
.io_out_2832(dataOut[2832]),
.io_out_2833(dataOut[2833]),
.io_out_2834(dataOut[2834]),
.io_out_2835(dataOut[2835]),
.io_out_2836(dataOut[2836]),
.io_out_2837(dataOut[2837]),
.io_out_2838(dataOut[2838]),
.io_out_2839(dataOut[2839]),
.io_out_2840(dataOut[2840]),
.io_out_2841(dataOut[2841]),
.io_out_2842(dataOut[2842]),
.io_out_2843(dataOut[2843]),
.io_out_2844(dataOut[2844]),
.io_out_2845(dataOut[2845]),
.io_out_2846(dataOut[2846]),
.io_out_2847(dataOut[2847]),
.io_out_2848(dataOut[2848]),
.io_out_2849(dataOut[2849]),
.io_out_2850(dataOut[2850]),
.io_out_2851(dataOut[2851]),
.io_out_2852(dataOut[2852]),
.io_out_2853(dataOut[2853]),
.io_out_2854(dataOut[2854]),
.io_out_2855(dataOut[2855]),
.io_out_2856(dataOut[2856]),
.io_out_2857(dataOut[2857]),
.io_out_2858(dataOut[2858]),
.io_out_2859(dataOut[2859]),
.io_out_2860(dataOut[2860]),
.io_out_2861(dataOut[2861]),
.io_out_2862(dataOut[2862]),
.io_out_2863(dataOut[2863]),
.io_out_2864(dataOut[2864]),
.io_out_2865(dataOut[2865]),
.io_out_2866(dataOut[2866]),
.io_out_2867(dataOut[2867]),
.io_out_2868(dataOut[2868]),
.io_out_2869(dataOut[2869]),
.io_out_2870(dataOut[2870]),
.io_out_2871(dataOut[2871]),
.io_out_2872(dataOut[2872]),
.io_out_2873(dataOut[2873]),
.io_out_2874(dataOut[2874]),
.io_out_2875(dataOut[2875]),
.io_out_2876(dataOut[2876]),
.io_out_2877(dataOut[2877]),
.io_out_2878(dataOut[2878]),
.io_out_2879(dataOut[2879]),
.io_out_2880(dataOut[2880]),
.io_out_2881(dataOut[2881]),
.io_out_2882(dataOut[2882]),
.io_out_2883(dataOut[2883]),
.io_out_2884(dataOut[2884]),
.io_out_2885(dataOut[2885]),
.io_out_2886(dataOut[2886]),
.io_out_2887(dataOut[2887]),
.io_out_2888(dataOut[2888]),
.io_out_2889(dataOut[2889]),
.io_out_2890(dataOut[2890]),
.io_out_2891(dataOut[2891]),
.io_out_2892(dataOut[2892]),
.io_out_2893(dataOut[2893]),
.io_out_2894(dataOut[2894]),
.io_out_2895(dataOut[2895]),
.io_out_2896(dataOut[2896]),
.io_out_2897(dataOut[2897]),
.io_out_2898(dataOut[2898]),
.io_out_2899(dataOut[2899]),
.io_out_2900(dataOut[2900]),
.io_out_2901(dataOut[2901]),
.io_out_2902(dataOut[2902]),
.io_out_2903(dataOut[2903]),
.io_out_2904(dataOut[2904]),
.io_out_2905(dataOut[2905]),
.io_out_2906(dataOut[2906]),
.io_out_2907(dataOut[2907]),
.io_out_2908(dataOut[2908]),
.io_out_2909(dataOut[2909]),
.io_out_2910(dataOut[2910]),
.io_out_2911(dataOut[2911]),
.io_out_2912(dataOut[2912]),
.io_out_2913(dataOut[2913]),
.io_out_2914(dataOut[2914]),
.io_out_2915(dataOut[2915]),
.io_out_2916(dataOut[2916]),
.io_out_2917(dataOut[2917]),
.io_out_2918(dataOut[2918]),
.io_out_2919(dataOut[2919]),
.io_out_2920(dataOut[2920]),
.io_out_2921(dataOut[2921]),
.io_out_2922(dataOut[2922]),
.io_out_2923(dataOut[2923]),
.io_out_2924(dataOut[2924]),
.io_out_2925(dataOut[2925]),
.io_out_2926(dataOut[2926]),
.io_out_2927(dataOut[2927]),
.io_out_2928(dataOut[2928]),
.io_out_2929(dataOut[2929]),
.io_out_2930(dataOut[2930]),
.io_out_2931(dataOut[2931]),
.io_out_2932(dataOut[2932]),
.io_out_2933(dataOut[2933]),
.io_out_2934(dataOut[2934]),
.io_out_2935(dataOut[2935]),
.io_out_2936(dataOut[2936]),
.io_out_2937(dataOut[2937]),
.io_out_2938(dataOut[2938]),
.io_out_2939(dataOut[2939]),
.io_out_2940(dataOut[2940]),
.io_out_2941(dataOut[2941]),
.io_out_2942(dataOut[2942]),
.io_out_2943(dataOut[2943]),
.io_out_2944(dataOut[2944]),
.io_out_2945(dataOut[2945]),
.io_out_2946(dataOut[2946]),
.io_out_2947(dataOut[2947]),
.io_out_2948(dataOut[2948]),
.io_out_2949(dataOut[2949]),
.io_out_2950(dataOut[2950]),
.io_out_2951(dataOut[2951]),
.io_out_2952(dataOut[2952]),
.io_out_2953(dataOut[2953]),
.io_out_2954(dataOut[2954]),
.io_out_2955(dataOut[2955]),
.io_out_2956(dataOut[2956]),
.io_out_2957(dataOut[2957]),
.io_out_2958(dataOut[2958]),
.io_out_2959(dataOut[2959]),
.io_out_2960(dataOut[2960]),
.io_out_2961(dataOut[2961]),
.io_out_2962(dataOut[2962]),
.io_out_2963(dataOut[2963]),
.io_out_2964(dataOut[2964]),
.io_out_2965(dataOut[2965]),
.io_out_2966(dataOut[2966]),
.io_out_2967(dataOut[2967]),
.io_out_2968(dataOut[2968]),
.io_out_2969(dataOut[2969]),
.io_out_2970(dataOut[2970]),
.io_out_2971(dataOut[2971]),
.io_out_2972(dataOut[2972]),
.io_out_2973(dataOut[2973]),
.io_out_2974(dataOut[2974]),
.io_out_2975(dataOut[2975]),
.io_out_2976(dataOut[2976]),
.io_out_2977(dataOut[2977]),
.io_out_2978(dataOut[2978]),
.io_out_2979(dataOut[2979]),
.io_out_2980(dataOut[2980]),
.io_out_2981(dataOut[2981]),
.io_out_2982(dataOut[2982]),
.io_out_2983(dataOut[2983]),
.io_out_2984(dataOut[2984]),
.io_out_2985(dataOut[2985]),
.io_out_2986(dataOut[2986]),
.io_out_2987(dataOut[2987]),
.io_out_2988(dataOut[2988]),
.io_out_2989(dataOut[2989]),
.io_out_2990(dataOut[2990]),
.io_out_2991(dataOut[2991]),
.io_out_2992(dataOut[2992]),
.io_out_2993(dataOut[2993]),
.io_out_2994(dataOut[2994]),
.io_out_2995(dataOut[2995]),
.io_out_2996(dataOut[2996]),
.io_out_2997(dataOut[2997]),
.io_out_2998(dataOut[2998]),
.io_out_2999(dataOut[2999]),
.io_out_3000(dataOut[3000]),
.io_out_3001(dataOut[3001]),
.io_out_3002(dataOut[3002]),
.io_out_3003(dataOut[3003]),
.io_out_3004(dataOut[3004]),
.io_out_3005(dataOut[3005]),
.io_out_3006(dataOut[3006]),
.io_out_3007(dataOut[3007]),
.io_out_3008(dataOut[3008]),
.io_out_3009(dataOut[3009]),
.io_out_3010(dataOut[3010]),
.io_out_3011(dataOut[3011]),
.io_out_3012(dataOut[3012]),
.io_out_3013(dataOut[3013]),
.io_out_3014(dataOut[3014]),
.io_out_3015(dataOut[3015]),
.io_out_3016(dataOut[3016]),
.io_out_3017(dataOut[3017]),
.io_out_3018(dataOut[3018]),
.io_out_3019(dataOut[3019]),
.io_out_3020(dataOut[3020]),
.io_out_3021(dataOut[3021]),
.io_out_3022(dataOut[3022]),
.io_out_3023(dataOut[3023]),
.io_out_3024(dataOut[3024]),
.io_out_3025(dataOut[3025]),
.io_out_3026(dataOut[3026]),
.io_out_3027(dataOut[3027]),
.io_out_3028(dataOut[3028]),
.io_out_3029(dataOut[3029]),
.io_out_3030(dataOut[3030]),
.io_out_3031(dataOut[3031]),
.io_out_3032(dataOut[3032]),
.io_out_3033(dataOut[3033]),
.io_out_3034(dataOut[3034]),
.io_out_3035(dataOut[3035]),
.io_out_3036(dataOut[3036]),
.io_out_3037(dataOut[3037]),
.io_out_3038(dataOut[3038]),
.io_out_3039(dataOut[3039]),
.io_out_3040(dataOut[3040]),
.io_out_3041(dataOut[3041]),
.io_out_3042(dataOut[3042]),
.io_out_3043(dataOut[3043]),
.io_out_3044(dataOut[3044]),
.io_out_3045(dataOut[3045]),
.io_out_3046(dataOut[3046]),
.io_out_3047(dataOut[3047]),
.io_out_3048(dataOut[3048]),
.io_out_3049(dataOut[3049]),
.io_out_3050(dataOut[3050]),
.io_out_3051(dataOut[3051]),
.io_out_3052(dataOut[3052]),
.io_out_3053(dataOut[3053]),
.io_out_3054(dataOut[3054]),
.io_out_3055(dataOut[3055]),
.io_out_3056(dataOut[3056]),
.io_out_3057(dataOut[3057]),
.io_out_3058(dataOut[3058]),
.io_out_3059(dataOut[3059]),
.io_out_3060(dataOut[3060]),
.io_out_3061(dataOut[3061]),
.io_out_3062(dataOut[3062]),
.io_out_3063(dataOut[3063]),
.io_out_3064(dataOut[3064]),
.io_out_3065(dataOut[3065]),
.io_out_3066(dataOut[3066]),
.io_out_3067(dataOut[3067]),
.io_out_3068(dataOut[3068]),
.io_out_3069(dataOut[3069]),
.io_out_3070(dataOut[3070]),
.io_out_3071(dataOut[3071]),
.io_out_3072(dataOut[3072]),
.io_out_3073(dataOut[3073]),
.io_out_3074(dataOut[3074]),
.io_out_3075(dataOut[3075]),
.io_out_3076(dataOut[3076]),
.io_out_3077(dataOut[3077]),
.io_out_3078(dataOut[3078]),
.io_out_3079(dataOut[3079]),
.io_out_3080(dataOut[3080]),
.io_out_3081(dataOut[3081]),
.io_out_3082(dataOut[3082]),
.io_out_3083(dataOut[3083]),
.io_out_3084(dataOut[3084]),
.io_out_3085(dataOut[3085]),
.io_out_3086(dataOut[3086]),
.io_out_3087(dataOut[3087]),
.io_out_3088(dataOut[3088]),
.io_out_3089(dataOut[3089]),
.io_out_3090(dataOut[3090]),
.io_out_3091(dataOut[3091]),
.io_out_3092(dataOut[3092]),
.io_out_3093(dataOut[3093]),
.io_out_3094(dataOut[3094]),
.io_out_3095(dataOut[3095]),
.io_out_3096(dataOut[3096]),
.io_out_3097(dataOut[3097]),
.io_out_3098(dataOut[3098]),
.io_out_3099(dataOut[3099]),
.io_out_3100(dataOut[3100]),
.io_out_3101(dataOut[3101]),
.io_out_3102(dataOut[3102]),
.io_out_3103(dataOut[3103]),
.io_out_3104(dataOut[3104]),
.io_out_3105(dataOut[3105]),
.io_out_3106(dataOut[3106]),
.io_out_3107(dataOut[3107]),
.io_out_3108(dataOut[3108]),
.io_out_3109(dataOut[3109]),
.io_out_3110(dataOut[3110]),
.io_out_3111(dataOut[3111]),
.io_out_3112(dataOut[3112]),
.io_out_3113(dataOut[3113]),
.io_out_3114(dataOut[3114]),
.io_out_3115(dataOut[3115]),
.io_out_3116(dataOut[3116]),
.io_out_3117(dataOut[3117]),
.io_out_3118(dataOut[3118]),
.io_out_3119(dataOut[3119]),
.io_out_3120(dataOut[3120]),
.io_out_3121(dataOut[3121]),
.io_out_3122(dataOut[3122]),
.io_out_3123(dataOut[3123]),
.io_out_3124(dataOut[3124]),
.io_out_3125(dataOut[3125]),
.io_out_3126(dataOut[3126]),
.io_out_3127(dataOut[3127]),
.io_out_3128(dataOut[3128]),
.io_out_3129(dataOut[3129]),
.io_out_3130(dataOut[3130]),
.io_out_3131(dataOut[3131]),
.io_out_3132(dataOut[3132]),
.io_out_3133(dataOut[3133]),
.io_out_3134(dataOut[3134]),
.io_out_3135(dataOut[3135]),
.io_out_3136(dataOut[3136]),
.io_out_3137(dataOut[3137]),
.io_out_3138(dataOut[3138]),
.io_out_3139(dataOut[3139]),
.io_out_3140(dataOut[3140]),
.io_out_3141(dataOut[3141]),
.io_out_3142(dataOut[3142]),
.io_out_3143(dataOut[3143]),
.io_out_3144(dataOut[3144]),
.io_out_3145(dataOut[3145]),
.io_out_3146(dataOut[3146]),
.io_out_3147(dataOut[3147]),
.io_out_3148(dataOut[3148]),
.io_out_3149(dataOut[3149]),
.io_out_3150(dataOut[3150]),
.io_out_3151(dataOut[3151]),
.io_out_3152(dataOut[3152]),
.io_out_3153(dataOut[3153]),
.io_out_3154(dataOut[3154]),
.io_out_3155(dataOut[3155]),
.io_out_3156(dataOut[3156]),
.io_out_3157(dataOut[3157]),
.io_out_3158(dataOut[3158]),
.io_out_3159(dataOut[3159]),
.io_out_3160(dataOut[3160]),
.io_out_3161(dataOut[3161]),
.io_out_3162(dataOut[3162]),
.io_out_3163(dataOut[3163]),
.io_out_3164(dataOut[3164]),
.io_out_3165(dataOut[3165]),
.io_out_3166(dataOut[3166]),
.io_out_3167(dataOut[3167]),
.io_out_3168(dataOut[3168]),
.io_out_3169(dataOut[3169]),
.io_out_3170(dataOut[3170]),
.io_out_3171(dataOut[3171]),
.io_out_3172(dataOut[3172]),
.io_out_3173(dataOut[3173]),
.io_out_3174(dataOut[3174]),
.io_out_3175(dataOut[3175]),
.io_out_3176(dataOut[3176]),
.io_out_3177(dataOut[3177]),
.io_out_3178(dataOut[3178]),
.io_out_3179(dataOut[3179]),
.io_out_3180(dataOut[3180]),
.io_out_3181(dataOut[3181]),
.io_out_3182(dataOut[3182]),
.io_out_3183(dataOut[3183]),
.io_out_3184(dataOut[3184]),
.io_out_3185(dataOut[3185]),
.io_out_3186(dataOut[3186]),
.io_out_3187(dataOut[3187]),
.io_out_3188(dataOut[3188]),
.io_out_3189(dataOut[3189]),
.io_out_3190(dataOut[3190]),
.io_out_3191(dataOut[3191]),
.io_out_3192(dataOut[3192]),
.io_out_3193(dataOut[3193]),
.io_out_3194(dataOut[3194]),
.io_out_3195(dataOut[3195]),
.io_out_3196(dataOut[3196]),
.io_out_3197(dataOut[3197]),
.io_out_3198(dataOut[3198]),
.io_out_3199(dataOut[3199]),
.io_out_3200(dataOut[3200]),
.io_out_3201(dataOut[3201]),
.io_out_3202(dataOut[3202]),
.io_out_3203(dataOut[3203]),
.io_out_3204(dataOut[3204]),
.io_out_3205(dataOut[3205]),
.io_out_3206(dataOut[3206]),
.io_out_3207(dataOut[3207]),
.io_out_3208(dataOut[3208]),
.io_out_3209(dataOut[3209]),
.io_out_3210(dataOut[3210]),
.io_out_3211(dataOut[3211]),
.io_out_3212(dataOut[3212]),
.io_out_3213(dataOut[3213]),
.io_out_3214(dataOut[3214]),
.io_out_3215(dataOut[3215]),
.io_out_3216(dataOut[3216]),
.io_out_3217(dataOut[3217]),
.io_out_3218(dataOut[3218]),
.io_out_3219(dataOut[3219]),
.io_out_3220(dataOut[3220]),
.io_out_3221(dataOut[3221]),
.io_out_3222(dataOut[3222]),
.io_out_3223(dataOut[3223]),
.io_out_3224(dataOut[3224]),
.io_out_3225(dataOut[3225]),
.io_out_3226(dataOut[3226]),
.io_out_3227(dataOut[3227]),
.io_out_3228(dataOut[3228]),
.io_out_3229(dataOut[3229]),
.io_out_3230(dataOut[3230]),
.io_out_3231(dataOut[3231]),
.io_out_3232(dataOut[3232]),
.io_out_3233(dataOut[3233]),
.io_out_3234(dataOut[3234]),
.io_out_3235(dataOut[3235]),
.io_out_3236(dataOut[3236]),
.io_out_3237(dataOut[3237]),
.io_out_3238(dataOut[3238]),
.io_out_3239(dataOut[3239]),
.io_out_3240(dataOut[3240]),
.io_out_3241(dataOut[3241]),
.io_out_3242(dataOut[3242]),
.io_out_3243(dataOut[3243]),
.io_out_3244(dataOut[3244]),
.io_out_3245(dataOut[3245]),
.io_out_3246(dataOut[3246]),
.io_out_3247(dataOut[3247]),
.io_out_3248(dataOut[3248]),
.io_out_3249(dataOut[3249]),
.io_out_3250(dataOut[3250]),
.io_out_3251(dataOut[3251]),
.io_out_3252(dataOut[3252]),
.io_out_3253(dataOut[3253]),
.io_out_3254(dataOut[3254]),
.io_out_3255(dataOut[3255]),
.io_out_3256(dataOut[3256]),
.io_out_3257(dataOut[3257]),
.io_out_3258(dataOut[3258]),
.io_out_3259(dataOut[3259]),
.io_out_3260(dataOut[3260]),
.io_out_3261(dataOut[3261]),
.io_out_3262(dataOut[3262]),
.io_out_3263(dataOut[3263]),
.io_out_3264(dataOut[3264]),
.io_out_3265(dataOut[3265]),
.io_out_3266(dataOut[3266]),
.io_out_3267(dataOut[3267]),
.io_out_3268(dataOut[3268]),
.io_out_3269(dataOut[3269]),
.io_out_3270(dataOut[3270]),
.io_out_3271(dataOut[3271]),
.io_out_3272(dataOut[3272]),
.io_out_3273(dataOut[3273]),
.io_out_3274(dataOut[3274]),
.io_out_3275(dataOut[3275]),
.io_out_3276(dataOut[3276]),
.io_out_3277(dataOut[3277]),
.io_out_3278(dataOut[3278]),
.io_out_3279(dataOut[3279]),
.io_out_3280(dataOut[3280]),
.io_out_3281(dataOut[3281]),
.io_out_3282(dataOut[3282]),
.io_out_3283(dataOut[3283]),
.io_out_3284(dataOut[3284]),
.io_out_3285(dataOut[3285]),
.io_out_3286(dataOut[3286]),
.io_out_3287(dataOut[3287]),
.io_out_3288(dataOut[3288]),
.io_out_3289(dataOut[3289]),
.io_out_3290(dataOut[3290]),
.io_out_3291(dataOut[3291]),
.io_out_3292(dataOut[3292]),
.io_out_3293(dataOut[3293]),
.io_out_3294(dataOut[3294]),
.io_out_3295(dataOut[3295]),
.io_out_3296(dataOut[3296]),
.io_out_3297(dataOut[3297]),
.io_out_3298(dataOut[3298]),
.io_out_3299(dataOut[3299]),
.io_out_3300(dataOut[3300]),
.io_out_3301(dataOut[3301]),
.io_out_3302(dataOut[3302]),
.io_out_3303(dataOut[3303]),
.io_out_3304(dataOut[3304]),
.io_out_3305(dataOut[3305]),
.io_out_3306(dataOut[3306]),
.io_out_3307(dataOut[3307]),
.io_out_3308(dataOut[3308]),
.io_out_3309(dataOut[3309]),
.io_out_3310(dataOut[3310]),
.io_out_3311(dataOut[3311]),
.io_out_3312(dataOut[3312]),
.io_out_3313(dataOut[3313]),
.io_out_3314(dataOut[3314]),
.io_out_3315(dataOut[3315]),
.io_out_3316(dataOut[3316]),
.io_out_3317(dataOut[3317]),
.io_out_3318(dataOut[3318]),
.io_out_3319(dataOut[3319]),
.io_out_3320(dataOut[3320]),
.io_out_3321(dataOut[3321]),
.io_out_3322(dataOut[3322]),
.io_out_3323(dataOut[3323]),
.io_out_3324(dataOut[3324]),
.io_out_3325(dataOut[3325]),
.io_out_3326(dataOut[3326]),
.io_out_3327(dataOut[3327]),
.io_out_3328(dataOut[3328]),
.io_out_3329(dataOut[3329]),
.io_out_3330(dataOut[3330]),
.io_out_3331(dataOut[3331]),
.io_out_3332(dataOut[3332]),
.io_out_3333(dataOut[3333]),
.io_out_3334(dataOut[3334]),
.io_out_3335(dataOut[3335]),
.io_out_3336(dataOut[3336]),
.io_out_3337(dataOut[3337]),
.io_out_3338(dataOut[3338]),
.io_out_3339(dataOut[3339]),
.io_out_3340(dataOut[3340]),
.io_out_3341(dataOut[3341]),
.io_out_3342(dataOut[3342]),
.io_out_3343(dataOut[3343]),
.io_out_3344(dataOut[3344]),
.io_out_3345(dataOut[3345]),
.io_out_3346(dataOut[3346]),
.io_out_3347(dataOut[3347]),
.io_out_3348(dataOut[3348]),
.io_out_3349(dataOut[3349]),
.io_out_3350(dataOut[3350]),
.io_out_3351(dataOut[3351]),
.io_out_3352(dataOut[3352]),
.io_out_3353(dataOut[3353]),
.io_out_3354(dataOut[3354]),
.io_out_3355(dataOut[3355]),
.io_out_3356(dataOut[3356]),
.io_out_3357(dataOut[3357]),
.io_out_3358(dataOut[3358]),
.io_out_3359(dataOut[3359]),
.io_out_3360(dataOut[3360]),
.io_out_3361(dataOut[3361]),
.io_out_3362(dataOut[3362]),
.io_out_3363(dataOut[3363]),
.io_out_3364(dataOut[3364]),
.io_out_3365(dataOut[3365]),
.io_out_3366(dataOut[3366]),
.io_out_3367(dataOut[3367]),
.io_out_3368(dataOut[3368]),
.io_out_3369(dataOut[3369]),
.io_out_3370(dataOut[3370]),
.io_out_3371(dataOut[3371]),
.io_out_3372(dataOut[3372]),
.io_out_3373(dataOut[3373]),
.io_out_3374(dataOut[3374]),
.io_out_3375(dataOut[3375]),
.io_out_3376(dataOut[3376]),
.io_out_3377(dataOut[3377]),
.io_out_3378(dataOut[3378]),
.io_out_3379(dataOut[3379]),
.io_out_3380(dataOut[3380]),
.io_out_3381(dataOut[3381]),
.io_out_3382(dataOut[3382]),
.io_out_3383(dataOut[3383]),
.io_out_3384(dataOut[3384]),
.io_out_3385(dataOut[3385]),
.io_out_3386(dataOut[3386]),
.io_out_3387(dataOut[3387]),
.io_out_3388(dataOut[3388]),
.io_out_3389(dataOut[3389]),
.io_out_3390(dataOut[3390]),
.io_out_3391(dataOut[3391]),
.io_out_3392(dataOut[3392]),
.io_out_3393(dataOut[3393]),
.io_out_3394(dataOut[3394]),
.io_out_3395(dataOut[3395]),
.io_out_3396(dataOut[3396]),
.io_out_3397(dataOut[3397]),
.io_out_3398(dataOut[3398]),
.io_out_3399(dataOut[3399]),
.io_out_3400(dataOut[3400]),
.io_out_3401(dataOut[3401]),
.io_out_3402(dataOut[3402]),
.io_out_3403(dataOut[3403]),
.io_out_3404(dataOut[3404]),
.io_out_3405(dataOut[3405]),
.io_out_3406(dataOut[3406]),
.io_out_3407(dataOut[3407]),
.io_out_3408(dataOut[3408]),
.io_out_3409(dataOut[3409]),
.io_out_3410(dataOut[3410]),
.io_out_3411(dataOut[3411]),
.io_out_3412(dataOut[3412]),
.io_out_3413(dataOut[3413]),
.io_out_3414(dataOut[3414]),
.io_out_3415(dataOut[3415]),
.io_out_3416(dataOut[3416]),
.io_out_3417(dataOut[3417]),
.io_out_3418(dataOut[3418]),
.io_out_3419(dataOut[3419]),
.io_out_3420(dataOut[3420]),
.io_out_3421(dataOut[3421]),
.io_out_3422(dataOut[3422]),
.io_out_3423(dataOut[3423]),
.io_out_3424(dataOut[3424]),
.io_out_3425(dataOut[3425]),
.io_out_3426(dataOut[3426]),
.io_out_3427(dataOut[3427]),
.io_out_3428(dataOut[3428]),
.io_out_3429(dataOut[3429]),
.io_out_3430(dataOut[3430]),
.io_out_3431(dataOut[3431]),
.io_out_3432(dataOut[3432]),
.io_out_3433(dataOut[3433]),
.io_out_3434(dataOut[3434]),
.io_out_3435(dataOut[3435]),
.io_out_3436(dataOut[3436]),
.io_out_3437(dataOut[3437]),
.io_out_3438(dataOut[3438]),
.io_out_3439(dataOut[3439]),
.io_out_3440(dataOut[3440]),
.io_out_3441(dataOut[3441]),
.io_out_3442(dataOut[3442]),
.io_out_3443(dataOut[3443]),
.io_out_3444(dataOut[3444]),
.io_out_3445(dataOut[3445]),
.io_out_3446(dataOut[3446]),
.io_out_3447(dataOut[3447]),
.io_out_3448(dataOut[3448]),
.io_out_3449(dataOut[3449]),
.io_out_3450(dataOut[3450]),
.io_out_3451(dataOut[3451]),
.io_out_3452(dataOut[3452]),
.io_out_3453(dataOut[3453]),
.io_out_3454(dataOut[3454]),
.io_out_3455(dataOut[3455]),
.io_out_3456(dataOut[3456]),
.io_out_3457(dataOut[3457]),
.io_out_3458(dataOut[3458]),
.io_out_3459(dataOut[3459]),
.io_out_3460(dataOut[3460]),
.io_out_3461(dataOut[3461]),
.io_out_3462(dataOut[3462]),
.io_out_3463(dataOut[3463]),
.io_out_3464(dataOut[3464]),
.io_out_3465(dataOut[3465]),
.io_out_3466(dataOut[3466]),
.io_out_3467(dataOut[3467]),
.io_out_3468(dataOut[3468]),
.io_out_3469(dataOut[3469]),
.io_out_3470(dataOut[3470]),
.io_out_3471(dataOut[3471]),
.io_out_3472(dataOut[3472]),
.io_out_3473(dataOut[3473]),
.io_out_3474(dataOut[3474]),
.io_out_3475(dataOut[3475]),
.io_out_3476(dataOut[3476]),
.io_out_3477(dataOut[3477]),
.io_out_3478(dataOut[3478]),
.io_out_3479(dataOut[3479]),
.io_out_3480(dataOut[3480]),
.io_out_3481(dataOut[3481]),
.io_out_3482(dataOut[3482]),
.io_out_3483(dataOut[3483]),
.io_out_3484(dataOut[3484]),
.io_out_3485(dataOut[3485]),
.io_out_3486(dataOut[3486]),
.io_out_3487(dataOut[3487]),
.io_out_3488(dataOut[3488]),
.io_out_3489(dataOut[3489]),
.io_out_3490(dataOut[3490]),
.io_out_3491(dataOut[3491]),
.io_out_3492(dataOut[3492]),
.io_out_3493(dataOut[3493]),
.io_out_3494(dataOut[3494]),
.io_out_3495(dataOut[3495]),
.io_out_3496(dataOut[3496]),
.io_out_3497(dataOut[3497]),
.io_out_3498(dataOut[3498]),
.io_out_3499(dataOut[3499]),
.io_out_3500(dataOut[3500]),
.io_out_3501(dataOut[3501]),
.io_out_3502(dataOut[3502]),
.io_out_3503(dataOut[3503]),
.io_out_3504(dataOut[3504]),
.io_out_3505(dataOut[3505]),
.io_out_3506(dataOut[3506]),
.io_out_3507(dataOut[3507]),
.io_out_3508(dataOut[3508]),
.io_out_3509(dataOut[3509]),
.io_out_3510(dataOut[3510]),
.io_out_3511(dataOut[3511]),
.io_out_3512(dataOut[3512]),
.io_out_3513(dataOut[3513]),
.io_out_3514(dataOut[3514]),
.io_out_3515(dataOut[3515]),
.io_out_3516(dataOut[3516]),
.io_out_3517(dataOut[3517]),
.io_out_3518(dataOut[3518]),
.io_out_3519(dataOut[3519]),
.io_out_3520(dataOut[3520]),
.io_out_3521(dataOut[3521]),
.io_out_3522(dataOut[3522]),
.io_out_3523(dataOut[3523]),
.io_out_3524(dataOut[3524]),
.io_out_3525(dataOut[3525]),
.io_out_3526(dataOut[3526]),
.io_out_3527(dataOut[3527]),
.io_out_3528(dataOut[3528]),
.io_out_3529(dataOut[3529]),
.io_out_3530(dataOut[3530]),
.io_out_3531(dataOut[3531]),
.io_out_3532(dataOut[3532]),
.io_out_3533(dataOut[3533]),
.io_out_3534(dataOut[3534]),
.io_out_3535(dataOut[3535]),
.io_out_3536(dataOut[3536]),
.io_out_3537(dataOut[3537]),
.io_out_3538(dataOut[3538]),
.io_out_3539(dataOut[3539]),
.io_out_3540(dataOut[3540]),
.io_out_3541(dataOut[3541]),
.io_out_3542(dataOut[3542]),
.io_out_3543(dataOut[3543]),
.io_out_3544(dataOut[3544]),
.io_out_3545(dataOut[3545]),
.io_out_3546(dataOut[3546]),
.io_out_3547(dataOut[3547]),
.io_out_3548(dataOut[3548]),
.io_out_3549(dataOut[3549]),
.io_out_3550(dataOut[3550]),
.io_out_3551(dataOut[3551]),
.io_out_3552(dataOut[3552]),
.io_out_3553(dataOut[3553]),
.io_out_3554(dataOut[3554]),
.io_out_3555(dataOut[3555]),
.io_out_3556(dataOut[3556]),
.io_out_3557(dataOut[3557]),
.io_out_3558(dataOut[3558]),
.io_out_3559(dataOut[3559]),
.io_out_3560(dataOut[3560]),
.io_out_3561(dataOut[3561]),
.io_out_3562(dataOut[3562]),
.io_out_3563(dataOut[3563]),
.io_out_3564(dataOut[3564]),
.io_out_3565(dataOut[3565]),
.io_out_3566(dataOut[3566]),
.io_out_3567(dataOut[3567]),
.io_out_3568(dataOut[3568]),
.io_out_3569(dataOut[3569]),
.io_out_3570(dataOut[3570]),
.io_out_3571(dataOut[3571]),
.io_out_3572(dataOut[3572]),
.io_out_3573(dataOut[3573]),
.io_out_3574(dataOut[3574]),
.io_out_3575(dataOut[3575]),
.io_out_3576(dataOut[3576]),
.io_out_3577(dataOut[3577]),
.io_out_3578(dataOut[3578]),
.io_out_3579(dataOut[3579]),
.io_out_3580(dataOut[3580]),
.io_out_3581(dataOut[3581]),
.io_out_3582(dataOut[3582]),
.io_out_3583(dataOut[3583]),
.io_out_3584(dataOut[3584]),
.io_out_3585(dataOut[3585]),
.io_out_3586(dataOut[3586]),
.io_out_3587(dataOut[3587]),
.io_out_3588(dataOut[3588]),
.io_out_3589(dataOut[3589]),
.io_out_3590(dataOut[3590]),
.io_out_3591(dataOut[3591]),
.io_out_3592(dataOut[3592]),
.io_out_3593(dataOut[3593]),
.io_out_3594(dataOut[3594]),
.io_out_3595(dataOut[3595]),
.io_out_3596(dataOut[3596]),
.io_out_3597(dataOut[3597]),
.io_out_3598(dataOut[3598]),
.io_out_3599(dataOut[3599]),
.io_out_3600(dataOut[3600]),
.io_out_3601(dataOut[3601]),
.io_out_3602(dataOut[3602]),
.io_out_3603(dataOut[3603]),
.io_out_3604(dataOut[3604]),
.io_out_3605(dataOut[3605]),
.io_out_3606(dataOut[3606]),
.io_out_3607(dataOut[3607]),
.io_out_3608(dataOut[3608]),
.io_out_3609(dataOut[3609]),
.io_out_3610(dataOut[3610]),
.io_out_3611(dataOut[3611]),
.io_out_3612(dataOut[3612]),
.io_out_3613(dataOut[3613]),
.io_out_3614(dataOut[3614]),
.io_out_3615(dataOut[3615]),
.io_out_3616(dataOut[3616]),
.io_out_3617(dataOut[3617]),
.io_out_3618(dataOut[3618]),
.io_out_3619(dataOut[3619]),
.io_out_3620(dataOut[3620]),
.io_out_3621(dataOut[3621]),
.io_out_3622(dataOut[3622]),
.io_out_3623(dataOut[3623]),
.io_out_3624(dataOut[3624]),
.io_out_3625(dataOut[3625]),
.io_out_3626(dataOut[3626]),
.io_out_3627(dataOut[3627]),
.io_out_3628(dataOut[3628]),
.io_out_3629(dataOut[3629]),
.io_out_3630(dataOut[3630]),
.io_out_3631(dataOut[3631]),
.io_out_3632(dataOut[3632]),
.io_out_3633(dataOut[3633]),
.io_out_3634(dataOut[3634]),
.io_out_3635(dataOut[3635]),
.io_out_3636(dataOut[3636]),
.io_out_3637(dataOut[3637]),
.io_out_3638(dataOut[3638]),
.io_out_3639(dataOut[3639]),
.io_out_3640(dataOut[3640]),
.io_out_3641(dataOut[3641]),
.io_out_3642(dataOut[3642]),
.io_out_3643(dataOut[3643]),
.io_out_3644(dataOut[3644]),
.io_out_3645(dataOut[3645]),
.io_out_3646(dataOut[3646]),
.io_out_3647(dataOut[3647]),
.io_out_3648(dataOut[3648]),
.io_out_3649(dataOut[3649]),
.io_out_3650(dataOut[3650]),
.io_out_3651(dataOut[3651]),
.io_out_3652(dataOut[3652]),
.io_out_3653(dataOut[3653]),
.io_out_3654(dataOut[3654]),
.io_out_3655(dataOut[3655]),
.io_out_3656(dataOut[3656]),
.io_out_3657(dataOut[3657]),
.io_out_3658(dataOut[3658]),
.io_out_3659(dataOut[3659]),
.io_out_3660(dataOut[3660]),
.io_out_3661(dataOut[3661]),
.io_out_3662(dataOut[3662]),
.io_out_3663(dataOut[3663]),
.io_out_3664(dataOut[3664]),
.io_out_3665(dataOut[3665]),
.io_out_3666(dataOut[3666]),
.io_out_3667(dataOut[3667]),
.io_out_3668(dataOut[3668]),
.io_out_3669(dataOut[3669]),
.io_out_3670(dataOut[3670]),
.io_out_3671(dataOut[3671]),
.io_out_3672(dataOut[3672]),
.io_out_3673(dataOut[3673]),
.io_out_3674(dataOut[3674]),
.io_out_3675(dataOut[3675]),
.io_out_3676(dataOut[3676]),
.io_out_3677(dataOut[3677]),
.io_out_3678(dataOut[3678]),
.io_out_3679(dataOut[3679]),
.io_out_3680(dataOut[3680]),
.io_out_3681(dataOut[3681]),
.io_out_3682(dataOut[3682]),
.io_out_3683(dataOut[3683]),
.io_out_3684(dataOut[3684]),
.io_out_3685(dataOut[3685]),
.io_out_3686(dataOut[3686]),
.io_out_3687(dataOut[3687]),
.io_out_3688(dataOut[3688]),
.io_out_3689(dataOut[3689]),
.io_out_3690(dataOut[3690]),
.io_out_3691(dataOut[3691]),
.io_out_3692(dataOut[3692]),
.io_out_3693(dataOut[3693]),
.io_out_3694(dataOut[3694]),
.io_out_3695(dataOut[3695]),
.io_out_3696(dataOut[3696]),
.io_out_3697(dataOut[3697]),
.io_out_3698(dataOut[3698]),
.io_out_3699(dataOut[3699]),
.io_out_3700(dataOut[3700]),
.io_out_3701(dataOut[3701]),
.io_out_3702(dataOut[3702]),
.io_out_3703(dataOut[3703]),
.io_out_3704(dataOut[3704]),
.io_out_3705(dataOut[3705]),
.io_out_3706(dataOut[3706]),
.io_out_3707(dataOut[3707]),
.io_out_3708(dataOut[3708]),
.io_out_3709(dataOut[3709]),
.io_out_3710(dataOut[3710]),
.io_out_3711(dataOut[3711]),
.io_out_3712(dataOut[3712]),
.io_out_3713(dataOut[3713]),
.io_out_3714(dataOut[3714]),
.io_out_3715(dataOut[3715]),
.io_out_3716(dataOut[3716]),
.io_out_3717(dataOut[3717]),
.io_out_3718(dataOut[3718]),
.io_out_3719(dataOut[3719]),
.io_out_3720(dataOut[3720]),
.io_out_3721(dataOut[3721]),
.io_out_3722(dataOut[3722]),
.io_out_3723(dataOut[3723]),
.io_out_3724(dataOut[3724]),
.io_out_3725(dataOut[3725]),
.io_out_3726(dataOut[3726]),
.io_out_3727(dataOut[3727]),
.io_out_3728(dataOut[3728]),
.io_out_3729(dataOut[3729]),
.io_out_3730(dataOut[3730]),
.io_out_3731(dataOut[3731]),
.io_out_3732(dataOut[3732]),
.io_out_3733(dataOut[3733]),
.io_out_3734(dataOut[3734]),
.io_out_3735(dataOut[3735]),
.io_out_3736(dataOut[3736]),
.io_out_3737(dataOut[3737]),
.io_out_3738(dataOut[3738]),
.io_out_3739(dataOut[3739]),
.io_out_3740(dataOut[3740]),
.io_out_3741(dataOut[3741]),
.io_out_3742(dataOut[3742]),
.io_out_3743(dataOut[3743]),
.io_out_3744(dataOut[3744]),
.io_out_3745(dataOut[3745]),
.io_out_3746(dataOut[3746]),
.io_out_3747(dataOut[3747]),
.io_out_3748(dataOut[3748]),
.io_out_3749(dataOut[3749]),
.io_out_3750(dataOut[3750]),
.io_out_3751(dataOut[3751]),
.io_out_3752(dataOut[3752]),
.io_out_3753(dataOut[3753]),
.io_out_3754(dataOut[3754]),
.io_out_3755(dataOut[3755]),
.io_out_3756(dataOut[3756]),
.io_out_3757(dataOut[3757]),
.io_out_3758(dataOut[3758]),
.io_out_3759(dataOut[3759]),
.io_out_3760(dataOut[3760]),
.io_out_3761(dataOut[3761]),
.io_out_3762(dataOut[3762]),
.io_out_3763(dataOut[3763]),
.io_out_3764(dataOut[3764]),
.io_out_3765(dataOut[3765]),
.io_out_3766(dataOut[3766]),
.io_out_3767(dataOut[3767]),
.io_out_3768(dataOut[3768]),
.io_out_3769(dataOut[3769]),
.io_out_3770(dataOut[3770]),
.io_out_3771(dataOut[3771]),
.io_out_3772(dataOut[3772]),
.io_out_3773(dataOut[3773]),
.io_out_3774(dataOut[3774]),
.io_out_3775(dataOut[3775]),
.io_out_3776(dataOut[3776]),
.io_out_3777(dataOut[3777]),
.io_out_3778(dataOut[3778]),
.io_out_3779(dataOut[3779]),
.io_out_3780(dataOut[3780]),
.io_out_3781(dataOut[3781]),
.io_out_3782(dataOut[3782]),
.io_out_3783(dataOut[3783]),
.io_out_3784(dataOut[3784]),
.io_out_3785(dataOut[3785]),
.io_out_3786(dataOut[3786]),
.io_out_3787(dataOut[3787]),
.io_out_3788(dataOut[3788]),
.io_out_3789(dataOut[3789]),
.io_out_3790(dataOut[3790]),
.io_out_3791(dataOut[3791]),
.io_out_3792(dataOut[3792]),
.io_out_3793(dataOut[3793]),
.io_out_3794(dataOut[3794]),
.io_out_3795(dataOut[3795]),
.io_out_3796(dataOut[3796]),
.io_out_3797(dataOut[3797]),
.io_out_3798(dataOut[3798]),
.io_out_3799(dataOut[3799]),
.io_out_3800(dataOut[3800]),
.io_out_3801(dataOut[3801]),
.io_out_3802(dataOut[3802]),
.io_out_3803(dataOut[3803]),
.io_out_3804(dataOut[3804]),
.io_out_3805(dataOut[3805]),
.io_out_3806(dataOut[3806]),
.io_out_3807(dataOut[3807]),
.io_out_3808(dataOut[3808]),
.io_out_3809(dataOut[3809]),
.io_out_3810(dataOut[3810]),
.io_out_3811(dataOut[3811]),
.io_out_3812(dataOut[3812]),
.io_out_3813(dataOut[3813]),
.io_out_3814(dataOut[3814]),
.io_out_3815(dataOut[3815]),
.io_out_3816(dataOut[3816]),
.io_out_3817(dataOut[3817]),
.io_out_3818(dataOut[3818]),
.io_out_3819(dataOut[3819]),
.io_out_3820(dataOut[3820]),
.io_out_3821(dataOut[3821]),
.io_out_3822(dataOut[3822]),
.io_out_3823(dataOut[3823]),
.io_out_3824(dataOut[3824]),
.io_out_3825(dataOut[3825]),
.io_out_3826(dataOut[3826]),
.io_out_3827(dataOut[3827]),
.io_out_3828(dataOut[3828]),
.io_out_3829(dataOut[3829]),
.io_out_3830(dataOut[3830]),
.io_out_3831(dataOut[3831]),
.io_out_3832(dataOut[3832]),
.io_out_3833(dataOut[3833]),
.io_out_3834(dataOut[3834]),
.io_out_3835(dataOut[3835]),
.io_out_3836(dataOut[3836]),
.io_out_3837(dataOut[3837]),
.io_out_3838(dataOut[3838]),
.io_out_3839(dataOut[3839]),
.io_out_3840(dataOut[3840]),
.io_out_3841(dataOut[3841]),
.io_out_3842(dataOut[3842]),
.io_out_3843(dataOut[3843]),
.io_out_3844(dataOut[3844]),
.io_out_3845(dataOut[3845]),
.io_out_3846(dataOut[3846]),
.io_out_3847(dataOut[3847]),
.io_out_3848(dataOut[3848]),
.io_out_3849(dataOut[3849]),
.io_out_3850(dataOut[3850]),
.io_out_3851(dataOut[3851]),
.io_out_3852(dataOut[3852]),
.io_out_3853(dataOut[3853]),
.io_out_3854(dataOut[3854]),
.io_out_3855(dataOut[3855]),
.io_out_3856(dataOut[3856]),
.io_out_3857(dataOut[3857]),
.io_out_3858(dataOut[3858]),
.io_out_3859(dataOut[3859]),
.io_out_3860(dataOut[3860]),
.io_out_3861(dataOut[3861]),
.io_out_3862(dataOut[3862]),
.io_out_3863(dataOut[3863]),
.io_out_3864(dataOut[3864]),
.io_out_3865(dataOut[3865]),
.io_out_3866(dataOut[3866]),
.io_out_3867(dataOut[3867]),
.io_out_3868(dataOut[3868]),
.io_out_3869(dataOut[3869]),
.io_out_3870(dataOut[3870]),
.io_out_3871(dataOut[3871]),
.io_out_3872(dataOut[3872]),
.io_out_3873(dataOut[3873]),
.io_out_3874(dataOut[3874]),
.io_out_3875(dataOut[3875]),
.io_out_3876(dataOut[3876]),
.io_out_3877(dataOut[3877]),
.io_out_3878(dataOut[3878]),
.io_out_3879(dataOut[3879]),
.io_out_3880(dataOut[3880]),
.io_out_3881(dataOut[3881]),
.io_out_3882(dataOut[3882]),
.io_out_3883(dataOut[3883]),
.io_out_3884(dataOut[3884]),
.io_out_3885(dataOut[3885]),
.io_out_3886(dataOut[3886]),
.io_out_3887(dataOut[3887]),
.io_out_3888(dataOut[3888]),
.io_out_3889(dataOut[3889]),
.io_out_3890(dataOut[3890]),
.io_out_3891(dataOut[3891]),
.io_out_3892(dataOut[3892]),
.io_out_3893(dataOut[3893]),
.io_out_3894(dataOut[3894]),
.io_out_3895(dataOut[3895]),
.io_out_3896(dataOut[3896]),
.io_out_3897(dataOut[3897]),
.io_out_3898(dataOut[3898]),
.io_out_3899(dataOut[3899]),
.io_out_3900(dataOut[3900]),
.io_out_3901(dataOut[3901]),
.io_out_3902(dataOut[3902]),
.io_out_3903(dataOut[3903]),
.io_out_3904(dataOut[3904]),
.io_out_3905(dataOut[3905]),
.io_out_3906(dataOut[3906]),
.io_out_3907(dataOut[3907]),
.io_out_3908(dataOut[3908]),
.io_out_3909(dataOut[3909]),
.io_out_3910(dataOut[3910]),
.io_out_3911(dataOut[3911]),
.io_out_3912(dataOut[3912]),
.io_out_3913(dataOut[3913]),
.io_out_3914(dataOut[3914]),
.io_out_3915(dataOut[3915]),
.io_out_3916(dataOut[3916]),
.io_out_3917(dataOut[3917]),
.io_out_3918(dataOut[3918]),
.io_out_3919(dataOut[3919]),
.io_out_3920(dataOut[3920]),
.io_out_3921(dataOut[3921]),
.io_out_3922(dataOut[3922]),
.io_out_3923(dataOut[3923]),
.io_out_3924(dataOut[3924]),
.io_out_3925(dataOut[3925]),
.io_out_3926(dataOut[3926]),
.io_out_3927(dataOut[3927]),
.io_out_3928(dataOut[3928]),
.io_out_3929(dataOut[3929]),
.io_out_3930(dataOut[3930]),
.io_out_3931(dataOut[3931]),
.io_out_3932(dataOut[3932]),
.io_out_3933(dataOut[3933]),
.io_out_3934(dataOut[3934]),
.io_out_3935(dataOut[3935]),
.io_out_3936(dataOut[3936]),
.io_out_3937(dataOut[3937]),
.io_out_3938(dataOut[3938]),
.io_out_3939(dataOut[3939]),
.io_out_3940(dataOut[3940]),
.io_out_3941(dataOut[3941]),
.io_out_3942(dataOut[3942]),
.io_out_3943(dataOut[3943]),
.io_out_3944(dataOut[3944]),
.io_out_3945(dataOut[3945]),
.io_out_3946(dataOut[3946]),
.io_out_3947(dataOut[3947]),
.io_out_3948(dataOut[3948]),
.io_out_3949(dataOut[3949]),
.io_out_3950(dataOut[3950]),
.io_out_3951(dataOut[3951]),
.io_out_3952(dataOut[3952]),
.io_out_3953(dataOut[3953]),
.io_out_3954(dataOut[3954]),
.io_out_3955(dataOut[3955]),
.io_out_3956(dataOut[3956]),
.io_out_3957(dataOut[3957]),
.io_out_3958(dataOut[3958]),
.io_out_3959(dataOut[3959]),
.io_out_3960(dataOut[3960]),
.io_out_3961(dataOut[3961]),
.io_out_3962(dataOut[3962]),
.io_out_3963(dataOut[3963]),
.io_out_3964(dataOut[3964]),
.io_out_3965(dataOut[3965]),
.io_out_3966(dataOut[3966]),
.io_out_3967(dataOut[3967]),
.io_out_3968(dataOut[3968]),
.io_out_3969(dataOut[3969]),
.io_out_3970(dataOut[3970]),
.io_out_3971(dataOut[3971]),
.io_out_3972(dataOut[3972]),
.io_out_3973(dataOut[3973]),
.io_out_3974(dataOut[3974]),
.io_out_3975(dataOut[3975]),
.io_out_3976(dataOut[3976]),
.io_out_3977(dataOut[3977]),
.io_out_3978(dataOut[3978]),
.io_out_3979(dataOut[3979]),
.io_out_3980(dataOut[3980]),
.io_out_3981(dataOut[3981]),
.io_out_3982(dataOut[3982]),
.io_out_3983(dataOut[3983]),
.io_out_3984(dataOut[3984]),
.io_out_3985(dataOut[3985]),
.io_out_3986(dataOut[3986]),
.io_out_3987(dataOut[3987]),
.io_out_3988(dataOut[3988]),
.io_out_3989(dataOut[3989]),
.io_out_3990(dataOut[3990]),
.io_out_3991(dataOut[3991]),
.io_out_3992(dataOut[3992]),
.io_out_3993(dataOut[3993]),
.io_out_3994(dataOut[3994]),
.io_out_3995(dataOut[3995]),
.io_out_3996(dataOut[3996]),
.io_out_3997(dataOut[3997]),
.io_out_3998(dataOut[3998]),
.io_out_3999(dataOut[3999]),
.io_out_4000(dataOut[4000]),
.io_out_4001(dataOut[4001]),
.io_out_4002(dataOut[4002]),
.io_out_4003(dataOut[4003]),
.io_out_4004(dataOut[4004]),
.io_out_4005(dataOut[4005]),
.io_out_4006(dataOut[4006]),
.io_out_4007(dataOut[4007]),
.io_out_4008(dataOut[4008]),
.io_out_4009(dataOut[4009]),
.io_out_4010(dataOut[4010]),
.io_out_4011(dataOut[4011]),
.io_out_4012(dataOut[4012]),
.io_out_4013(dataOut[4013]),
.io_out_4014(dataOut[4014]),
.io_out_4015(dataOut[4015]),
.io_out_4016(dataOut[4016]),
.io_out_4017(dataOut[4017]),
.io_out_4018(dataOut[4018]),
.io_out_4019(dataOut[4019]),
.io_out_4020(dataOut[4020]),
.io_out_4021(dataOut[4021]),
.io_out_4022(dataOut[4022]),
.io_out_4023(dataOut[4023]),
.io_out_4024(dataOut[4024]),
.io_out_4025(dataOut[4025]),
.io_out_4026(dataOut[4026]),
.io_out_4027(dataOut[4027]),
.io_out_4028(dataOut[4028]),
.io_out_4029(dataOut[4029]),
.io_out_4030(dataOut[4030]),
.io_out_4031(dataOut[4031]),
.io_out_4032(dataOut[4032]),
.io_out_4033(dataOut[4033]),
.io_out_4034(dataOut[4034]),
.io_out_4035(dataOut[4035]),
.io_out_4036(dataOut[4036]),
.io_out_4037(dataOut[4037]),
.io_out_4038(dataOut[4038]),
.io_out_4039(dataOut[4039]),
.io_out_4040(dataOut[4040]),
.io_out_4041(dataOut[4041]),
.io_out_4042(dataOut[4042]),
.io_out_4043(dataOut[4043]),
.io_out_4044(dataOut[4044]),
.io_out_4045(dataOut[4045]),
.io_out_4046(dataOut[4046]),
.io_out_4047(dataOut[4047]),
.io_out_4048(dataOut[4048]),
.io_out_4049(dataOut[4049]),
.io_out_4050(dataOut[4050]),
.io_out_4051(dataOut[4051]),
.io_out_4052(dataOut[4052]),
.io_out_4053(dataOut[4053]),
.io_out_4054(dataOut[4054]),
.io_out_4055(dataOut[4055]),
.io_out_4056(dataOut[4056]),
.io_out_4057(dataOut[4057]),
.io_out_4058(dataOut[4058]),
.io_out_4059(dataOut[4059]),
.io_out_4060(dataOut[4060]),
.io_out_4061(dataOut[4061]),
.io_out_4062(dataOut[4062]),
.io_out_4063(dataOut[4063]),
.io_out_4064(dataOut[4064]),
.io_out_4065(dataOut[4065]),
.io_out_4066(dataOut[4066]),
.io_out_4067(dataOut[4067]),
.io_out_4068(dataOut[4068]),
.io_out_4069(dataOut[4069]),
.io_out_4070(dataOut[4070]),
.io_out_4071(dataOut[4071]),
.io_out_4072(dataOut[4072]),
.io_out_4073(dataOut[4073]),
.io_out_4074(dataOut[4074]),
.io_out_4075(dataOut[4075]),
.io_out_4076(dataOut[4076]),
.io_out_4077(dataOut[4077]),
.io_out_4078(dataOut[4078]),
.io_out_4079(dataOut[4079]),
.io_out_4080(dataOut[4080]),
.io_out_4081(dataOut[4081]),
.io_out_4082(dataOut[4082]),
.io_out_4083(dataOut[4083]),
.io_out_4084(dataOut[4084]),
.io_out_4085(dataOut[4085]),
.io_out_4086(dataOut[4086]),
.io_out_4087(dataOut[4087]),
.io_out_4088(dataOut[4088]),
.io_out_4089(dataOut[4089]),
.io_out_4090(dataOut[4090]),
.io_out_4091(dataOut[4091]),
.io_out_4092(dataOut[4092]),
.io_out_4093(dataOut[4093]),
.io_out_4094(dataOut[4094]),
.io_out_4095(dataOut[4095]),
.io_matchingBytes_0(matchingBytes[0]),
.io_matchingBytes_1(matchingBytes[1]),
.io_matchingBytes_2(matchingBytes[2]),
.io_matchingBytes_3(matchingBytes[3]),
.io_matchingBytes_4(matchingBytes[4]),
.io_matchingBytes_5(matchingBytes[5]),
.io_matchingBytes_6(matchingBytes[6]),
.io_matchingBytes_7(matchingBytes[7]),
.io_matchingBytes_8(matchingBytes[8]),
.io_matchingBytes_9(matchingBytes[9]),
.io_matchingBytes_10(matchingBytes[10]),
.io_matchingBytes_11(matchingBytes[11]),
.io_matchingBytes_12(matchingBytes[12]),
.io_matchingBytes_13(matchingBytes[13]),
.io_matchingBytes_14(matchingBytes[14]),
.io_matchingBytes_15(matchingBytes[15]),
.io_matchingBytes_16(matchingBytes[16]),
.io_matchingBytes_17(matchingBytes[17]),
.io_matchingBytes_18(matchingBytes[18]),
.io_matchingBytes_19(matchingBytes[19]),
.io_matchingBytes_20(matchingBytes[20]),
.io_matchingBytes_21(matchingBytes[21]),
.io_matchingBytes_22(matchingBytes[22]),
.io_matchingBytes_23(matchingBytes[23]),
.io_matchingBytes_24(matchingBytes[24]),
.io_matchingBytes_25(matchingBytes[25]),
.io_matchingBytes_26(matchingBytes[26]),
.io_matchingBytes_27(matchingBytes[27]),
.io_matchingBytes_28(matchingBytes[28]),
.io_matchingBytes_29(matchingBytes[29]),
.io_matchingBytes_30(matchingBytes[30]),
.io_matchingBytes_31(matchingBytes[31]),
.io_matchingBytes_32(matchingBytes[32]),
.io_matchingBytes_33(matchingBytes[33]),
.io_matchingBytes_34(matchingBytes[34]),
.io_matchingBytes_35(matchingBytes[35]),
.io_matchingBytes_36(matchingBytes[36]),
.io_matchingBytes_37(matchingBytes[37]),
.io_matchingBytes_38(matchingBytes[38]),
.io_matchingBytes_39(matchingBytes[39]),
.io_matchingBytes_40(matchingBytes[40]),
.io_matchingBytes_41(matchingBytes[41]),
.io_matchingBytes_42(matchingBytes[42]),
.io_matchingBytes_43(matchingBytes[43]),
.io_matchingBytes_44(matchingBytes[44]),
.io_matchingBytes_45(matchingBytes[45]),
.io_matchingBytes_46(matchingBytes[46]),
.io_matchingBytes_47(matchingBytes[47]),
.io_matchingBytes_48(matchingBytes[48]),
.io_matchingBytes_49(matchingBytes[49]),
.io_matchingBytes_50(matchingBytes[50]),
.io_matchingBytes_51(matchingBytes[51]),
.io_matchingBytes_52(matchingBytes[52]),
.io_matchingBytes_53(matchingBytes[53]),
.io_matchingBytes_54(matchingBytes[54]),
.io_matchingBytes_55(matchingBytes[55]),
.io_matchingBytes_56(matchingBytes[56]),
.io_matchingBytes_57(matchingBytes[57]),
.io_matchingBytes_58(matchingBytes[58]),
.io_matchingBytes_59(matchingBytes[59]),
.io_matchingBytes_60(matchingBytes[60]),
.io_matchingBytes_61(matchingBytes[61]),
.io_matchingBytes_62(matchingBytes[62]),
.io_matchingBytes_63(matchingBytes[63]),
.io_matchingBytes_64(matchingBytes[64]),
.io_matchingBytes_65(matchingBytes[65]),
.io_matchingBytes_66(matchingBytes[66]),
.io_matchingBytes_67(matchingBytes[67]),
.io_matchingBytes_68(matchingBytes[68]),
.io_matchingBytes_69(matchingBytes[69]),
.io_matchingBytes_70(matchingBytes[70]),
.io_matchingBytes_71(matchingBytes[71]),
.io_matchingBytes_72(matchingBytes[72]),
.io_matchingBytes_73(matchingBytes[73]),
.io_matchingBytes_74(matchingBytes[74]),
.io_matchingBytes_75(matchingBytes[75]),
.io_matchingBytes_76(matchingBytes[76]),
.io_matchingBytes_77(matchingBytes[77]),
.io_matchingBytes_78(matchingBytes[78]),
.io_matchingBytes_79(matchingBytes[79]),
.io_matchingBytes_80(matchingBytes[80]),
.io_matchingBytes_81(matchingBytes[81]),
.io_matchingBytes_82(matchingBytes[82]),
.io_matchingBytes_83(matchingBytes[83]),
.io_matchingBytes_84(matchingBytes[84]),
.io_matchingBytes_85(matchingBytes[85]),
.io_matchingBytes_86(matchingBytes[86]),
.io_matchingBytes_87(matchingBytes[87]),
.io_matchingBytes_88(matchingBytes[88]),
.io_matchingBytes_89(matchingBytes[89]),
.io_matchingBytes_90(matchingBytes[90]),
.io_matchingBytes_91(matchingBytes[91]),
.io_matchingBytes_92(matchingBytes[92]),
.io_matchingBytes_93(matchingBytes[93]),
.io_matchingBytes_94(matchingBytes[94]),
.io_matchingBytes_95(matchingBytes[95]),
.io_matchingBytes_96(matchingBytes[96]),
.io_matchingBytes_97(matchingBytes[97]),
.io_matchingBytes_98(matchingBytes[98]),
.io_matchingBytes_99(matchingBytes[99]),
.io_matchingBytes_100(matchingBytes[100]),
.io_matchingBytes_101(matchingBytes[101]),
.io_matchingBytes_102(matchingBytes[102]),
.io_matchingBytes_103(matchingBytes[103]),
.io_matchingBytes_104(matchingBytes[104]),
.io_matchingBytes_105(matchingBytes[105]),
.io_matchingBytes_106(matchingBytes[106]),
.io_matchingBytes_107(matchingBytes[107]),
.io_matchingBytes_108(matchingBytes[108]),
.io_matchingBytes_109(matchingBytes[109]),
.io_matchingBytes_110(matchingBytes[110]),
.io_matchingBytes_111(matchingBytes[111]),
.io_matchingBytes_112(matchingBytes[112]),
.io_matchingBytes_113(matchingBytes[113]),
.io_matchingBytes_114(matchingBytes[114]),
.io_matchingBytes_115(matchingBytes[115]),
.io_matchingBytes_116(matchingBytes[116]),
.io_matchingBytes_117(matchingBytes[117]),
.io_matchingBytes_118(matchingBytes[118]),
.io_matchingBytes_119(matchingBytes[119]),
.io_matchingBytes_120(matchingBytes[120]),
.io_matchingBytes_121(matchingBytes[121]),
.io_matchingBytes_122(matchingBytes[122]),
.io_matchingBytes_123(matchingBytes[123]),
.io_matchingBytes_124(matchingBytes[124]),
.io_matchingBytes_125(matchingBytes[125]),
.io_matchingBytes_126(matchingBytes[126]),
.io_matchingBytes_127(matchingBytes[127]),
.io_matchingBytes_128(matchingBytes[128]),
.io_matchingBytes_129(matchingBytes[129]),
.io_matchingBytes_130(matchingBytes[130]),
.io_matchingBytes_131(matchingBytes[131]),
.io_matchingBytes_132(matchingBytes[132]),
.io_matchingBytes_133(matchingBytes[133]),
.io_matchingBytes_134(matchingBytes[134]),
.io_matchingBytes_135(matchingBytes[135]),
.io_matchingBytes_136(matchingBytes[136]),
.io_matchingBytes_137(matchingBytes[137]),
.io_matchingBytes_138(matchingBytes[138]),
.io_matchingBytes_139(matchingBytes[139]),
.io_matchingBytes_140(matchingBytes[140]),
.io_matchingBytes_141(matchingBytes[141]),
.io_matchingBytes_142(matchingBytes[142]),
.io_matchingBytes_143(matchingBytes[143]),
.io_matchingBytes_144(matchingBytes[144]),
.io_matchingBytes_145(matchingBytes[145]),
.io_matchingBytes_146(matchingBytes[146]),
.io_matchingBytes_147(matchingBytes[147]),
.io_matchingBytes_148(matchingBytes[148]),
.io_matchingBytes_149(matchingBytes[149]),
.io_matchingBytes_150(matchingBytes[150]),
.io_matchingBytes_151(matchingBytes[151]),
.io_matchingBytes_152(matchingBytes[152]),
.io_matchingBytes_153(matchingBytes[153]),
.io_matchingBytes_154(matchingBytes[154]),
.io_matchingBytes_155(matchingBytes[155]),
.io_matchingBytes_156(matchingBytes[156]),
.io_matchingBytes_157(matchingBytes[157]),
.io_matchingBytes_158(matchingBytes[158]),
.io_matchingBytes_159(matchingBytes[159]),
.io_matchingBytes_160(matchingBytes[160]),
.io_matchingBytes_161(matchingBytes[161]),
.io_matchingBytes_162(matchingBytes[162]),
.io_matchingBytes_163(matchingBytes[163]),
.io_matchingBytes_164(matchingBytes[164]),
.io_matchingBytes_165(matchingBytes[165]),
.io_matchingBytes_166(matchingBytes[166]),
.io_matchingBytes_167(matchingBytes[167]),
.io_matchingBytes_168(matchingBytes[168]),
.io_matchingBytes_169(matchingBytes[169]),
.io_matchingBytes_170(matchingBytes[170]),
.io_matchingBytes_171(matchingBytes[171]),
.io_matchingBytes_172(matchingBytes[172]),
.io_matchingBytes_173(matchingBytes[173]),
.io_matchingBytes_174(matchingBytes[174]),
.io_matchingBytes_175(matchingBytes[175]),
.io_matchingBytes_176(matchingBytes[176]),
.io_matchingBytes_177(matchingBytes[177]),
.io_matchingBytes_178(matchingBytes[178]),
.io_matchingBytes_179(matchingBytes[179]),
.io_matchingBytes_180(matchingBytes[180]),
.io_matchingBytes_181(matchingBytes[181]),
.io_matchingBytes_182(matchingBytes[182]),
.io_matchingBytes_183(matchingBytes[183]),
.io_matchingBytes_184(matchingBytes[184]),
.io_matchingBytes_185(matchingBytes[185]),
.io_matchingBytes_186(matchingBytes[186]),
.io_matchingBytes_187(matchingBytes[187]),
.io_matchingBytes_188(matchingBytes[188]),
.io_matchingBytes_189(matchingBytes[189]),
.io_matchingBytes_190(matchingBytes[190]),
.io_matchingBytes_191(matchingBytes[191]),
.io_matchingBytes_192(matchingBytes[192]),
.io_matchingBytes_193(matchingBytes[193]),
.io_matchingBytes_194(matchingBytes[194]),
.io_matchingBytes_195(matchingBytes[195]),
.io_matchingBytes_196(matchingBytes[196]),
.io_matchingBytes_197(matchingBytes[197]),
.io_matchingBytes_198(matchingBytes[198]),
.io_matchingBytes_199(matchingBytes[199]),
.io_matchingBytes_200(matchingBytes[200]),
.io_matchingBytes_201(matchingBytes[201]),
.io_matchingBytes_202(matchingBytes[202]),
.io_matchingBytes_203(matchingBytes[203]),
.io_matchingBytes_204(matchingBytes[204]),
.io_matchingBytes_205(matchingBytes[205]),
.io_matchingBytes_206(matchingBytes[206]),
.io_matchingBytes_207(matchingBytes[207]),
.io_matchingBytes_208(matchingBytes[208]),
.io_matchingBytes_209(matchingBytes[209]),
.io_matchingBytes_210(matchingBytes[210]),
.io_matchingBytes_211(matchingBytes[211]),
.io_matchingBytes_212(matchingBytes[212]),
.io_matchingBytes_213(matchingBytes[213]),
.io_matchingBytes_214(matchingBytes[214]),
.io_matchingBytes_215(matchingBytes[215]),
.io_matchingBytes_216(matchingBytes[216]),
.io_matchingBytes_217(matchingBytes[217]),
.io_matchingBytes_218(matchingBytes[218]),
.io_matchingBytes_219(matchingBytes[219]),
.io_matchingBytes_220(matchingBytes[220]),
.io_matchingBytes_221(matchingBytes[221]),
.io_matchingBytes_222(matchingBytes[222]),
.io_matchingBytes_223(matchingBytes[223]),
.io_matchingBytes_224(matchingBytes[224]),
.io_matchingBytes_225(matchingBytes[225]),
.io_matchingBytes_226(matchingBytes[226]),
.io_matchingBytes_227(matchingBytes[227]),
.io_matchingBytes_228(matchingBytes[228]),
.io_matchingBytes_229(matchingBytes[229]),
.io_matchingBytes_230(matchingBytes[230]),
.io_matchingBytes_231(matchingBytes[231]),
.io_matchingBytes_232(matchingBytes[232]),
.io_matchingBytes_233(matchingBytes[233]),
.io_matchingBytes_234(matchingBytes[234]),
.io_matchingBytes_235(matchingBytes[235]),
.io_matchingBytes_236(matchingBytes[236]),
.io_matchingBytes_237(matchingBytes[237]),
.io_matchingBytes_238(matchingBytes[238]),
.io_matchingBytes_239(matchingBytes[239]),
.io_matchingBytes_240(matchingBytes[240]),
.io_matchingBytes_241(matchingBytes[241]),
.io_matchingBytes_242(matchingBytes[242]),
.io_matchingBytes_243(matchingBytes[243]),
.io_matchingBytes_244(matchingBytes[244]),
.io_matchingBytes_245(matchingBytes[245]),
.io_matchingBytes_246(matchingBytes[246]),
.io_matchingBytes_247(matchingBytes[247]),
.io_matchingBytes_248(matchingBytes[248]),
.io_matchingBytes_249(matchingBytes[249]),
.io_matchingBytes_250(matchingBytes[250]),
.io_matchingBytes_251(matchingBytes[251]),
.io_matchingBytes_252(matchingBytes[252]),
.io_matchingBytes_253(matchingBytes[253]),
.io_matchingBytes_254(matchingBytes[254]),
.io_matchingBytes_255(matchingBytes[255]),
.io_matchingBytes_256(matchingBytes[256]),
.io_matchingBytes_257(matchingBytes[257]),
.io_matchingBytes_258(matchingBytes[258]),
.io_matchingBytes_259(matchingBytes[259]),
.io_matchingBytes_260(matchingBytes[260]),
.io_matchingBytes_261(matchingBytes[261]),
.io_matchingBytes_262(matchingBytes[262]),
.io_matchingBytes_263(matchingBytes[263]),
.io_matchingBytes_264(matchingBytes[264]),
.io_matchingBytes_265(matchingBytes[265]),
.io_matchingBytes_266(matchingBytes[266]),
.io_matchingBytes_267(matchingBytes[267]),
.io_matchingBytes_268(matchingBytes[268]),
.io_matchingBytes_269(matchingBytes[269]),
.io_matchingBytes_270(matchingBytes[270]),
.io_matchingBytes_271(matchingBytes[271]),
.io_matchingBytes_272(matchingBytes[272]),
.io_matchingBytes_273(matchingBytes[273]),
.io_matchingBytes_274(matchingBytes[274]),
.io_matchingBytes_275(matchingBytes[275]),
.io_matchingBytes_276(matchingBytes[276]),
.io_matchingBytes_277(matchingBytes[277]),
.io_matchingBytes_278(matchingBytes[278]),
.io_matchingBytes_279(matchingBytes[279]),
.io_matchingBytes_280(matchingBytes[280]),
.io_matchingBytes_281(matchingBytes[281]),
.io_matchingBytes_282(matchingBytes[282]),
.io_matchingBytes_283(matchingBytes[283]),
.io_matchingBytes_284(matchingBytes[284]),
.io_matchingBytes_285(matchingBytes[285]),
.io_matchingBytes_286(matchingBytes[286]),
.io_matchingBytes_287(matchingBytes[287]),
.io_matchingBytes_288(matchingBytes[288]),
.io_matchingBytes_289(matchingBytes[289]),
.io_matchingBytes_290(matchingBytes[290]),
.io_matchingBytes_291(matchingBytes[291]),
.io_matchingBytes_292(matchingBytes[292]),
.io_matchingBytes_293(matchingBytes[293]),
.io_matchingBytes_294(matchingBytes[294]),
.io_matchingBytes_295(matchingBytes[295]),
.io_matchingBytes_296(matchingBytes[296]),
.io_matchingBytes_297(matchingBytes[297]),
.io_matchingBytes_298(matchingBytes[298]),
.io_matchingBytes_299(matchingBytes[299]),
.io_matchingBytes_300(matchingBytes[300]),
.io_matchingBytes_301(matchingBytes[301]),
.io_matchingBytes_302(matchingBytes[302]),
.io_matchingBytes_303(matchingBytes[303]),
.io_matchingBytes_304(matchingBytes[304]),
.io_matchingBytes_305(matchingBytes[305]),
.io_matchingBytes_306(matchingBytes[306]),
.io_matchingBytes_307(matchingBytes[307]),
.io_matchingBytes_308(matchingBytes[308]),
.io_matchingBytes_309(matchingBytes[309]),
.io_matchingBytes_310(matchingBytes[310]),
.io_matchingBytes_311(matchingBytes[311]),
.io_matchingBytes_312(matchingBytes[312]),
.io_matchingBytes_313(matchingBytes[313]),
.io_matchingBytes_314(matchingBytes[314]),
.io_matchingBytes_315(matchingBytes[315]),
.io_matchingBytes_316(matchingBytes[316]),
.io_matchingBytes_317(matchingBytes[317]),
.io_matchingBytes_318(matchingBytes[318]),
.io_matchingBytes_319(matchingBytes[319]),
.io_matchingBytes_320(matchingBytes[320]),
.io_matchingBytes_321(matchingBytes[321]),
.io_matchingBytes_322(matchingBytes[322]),
.io_matchingBytes_323(matchingBytes[323]),
.io_matchingBytes_324(matchingBytes[324]),
.io_matchingBytes_325(matchingBytes[325]),
.io_matchingBytes_326(matchingBytes[326]),
.io_matchingBytes_327(matchingBytes[327]),
.io_matchingBytes_328(matchingBytes[328]),
.io_matchingBytes_329(matchingBytes[329]),
.io_matchingBytes_330(matchingBytes[330]),
.io_matchingBytes_331(matchingBytes[331]),
.io_matchingBytes_332(matchingBytes[332]),
.io_matchingBytes_333(matchingBytes[333]),
.io_matchingBytes_334(matchingBytes[334]),
.io_matchingBytes_335(matchingBytes[335]),
.io_matchingBytes_336(matchingBytes[336]),
.io_matchingBytes_337(matchingBytes[337]),
.io_matchingBytes_338(matchingBytes[338]),
.io_matchingBytes_339(matchingBytes[339]),
.io_matchingBytes_340(matchingBytes[340]),
.io_matchingBytes_341(matchingBytes[341]),
.io_matchingBytes_342(matchingBytes[342]),
.io_matchingBytes_343(matchingBytes[343]),
.io_matchingBytes_344(matchingBytes[344]),
.io_matchingBytes_345(matchingBytes[345]),
.io_matchingBytes_346(matchingBytes[346]),
.io_matchingBytes_347(matchingBytes[347]),
.io_matchingBytes_348(matchingBytes[348]),
.io_matchingBytes_349(matchingBytes[349]),
.io_matchingBytes_350(matchingBytes[350]),
.io_matchingBytes_351(matchingBytes[351]),
.io_matchingBytes_352(matchingBytes[352]),
.io_matchingBytes_353(matchingBytes[353]),
.io_matchingBytes_354(matchingBytes[354]),
.io_matchingBytes_355(matchingBytes[355]),
.io_matchingBytes_356(matchingBytes[356]),
.io_matchingBytes_357(matchingBytes[357]),
.io_matchingBytes_358(matchingBytes[358]),
.io_matchingBytes_359(matchingBytes[359]),
.io_matchingBytes_360(matchingBytes[360]),
.io_matchingBytes_361(matchingBytes[361]),
.io_matchingBytes_362(matchingBytes[362]),
.io_matchingBytes_363(matchingBytes[363]),
.io_matchingBytes_364(matchingBytes[364]),
.io_matchingBytes_365(matchingBytes[365]),
.io_matchingBytes_366(matchingBytes[366]),
.io_matchingBytes_367(matchingBytes[367]),
.io_matchingBytes_368(matchingBytes[368]),
.io_matchingBytes_369(matchingBytes[369]),
.io_matchingBytes_370(matchingBytes[370]),
.io_matchingBytes_371(matchingBytes[371]),
.io_matchingBytes_372(matchingBytes[372]),
.io_matchingBytes_373(matchingBytes[373]),
.io_matchingBytes_374(matchingBytes[374]),
.io_matchingBytes_375(matchingBytes[375]),
.io_matchingBytes_376(matchingBytes[376]),
.io_matchingBytes_377(matchingBytes[377]),
.io_matchingBytes_378(matchingBytes[378]),
.io_matchingBytes_379(matchingBytes[379]),
.io_matchingBytes_380(matchingBytes[380]),
.io_matchingBytes_381(matchingBytes[381]),
.io_matchingBytes_382(matchingBytes[382]),
.io_matchingBytes_383(matchingBytes[383]),
.io_matchingBytes_384(matchingBytes[384]),
.io_matchingBytes_385(matchingBytes[385]),
.io_matchingBytes_386(matchingBytes[386]),
.io_matchingBytes_387(matchingBytes[387]),
.io_matchingBytes_388(matchingBytes[388]),
.io_matchingBytes_389(matchingBytes[389]),
.io_matchingBytes_390(matchingBytes[390]),
.io_matchingBytes_391(matchingBytes[391]),
.io_matchingBytes_392(matchingBytes[392]),
.io_matchingBytes_393(matchingBytes[393]),
.io_matchingBytes_394(matchingBytes[394]),
.io_matchingBytes_395(matchingBytes[395]),
.io_matchingBytes_396(matchingBytes[396]),
.io_matchingBytes_397(matchingBytes[397]),
.io_matchingBytes_398(matchingBytes[398]),
.io_matchingBytes_399(matchingBytes[399]),
.io_matchingBytes_400(matchingBytes[400]),
.io_matchingBytes_401(matchingBytes[401]),
.io_matchingBytes_402(matchingBytes[402]),
.io_matchingBytes_403(matchingBytes[403]),
.io_matchingBytes_404(matchingBytes[404]),
.io_matchingBytes_405(matchingBytes[405]),
.io_matchingBytes_406(matchingBytes[406]),
.io_matchingBytes_407(matchingBytes[407]),
.io_matchingBytes_408(matchingBytes[408]),
.io_matchingBytes_409(matchingBytes[409]),
.io_matchingBytes_410(matchingBytes[410]),
.io_matchingBytes_411(matchingBytes[411]),
.io_matchingBytes_412(matchingBytes[412]),
.io_matchingBytes_413(matchingBytes[413]),
.io_matchingBytes_414(matchingBytes[414]),
.io_matchingBytes_415(matchingBytes[415]),
.io_matchingBytes_416(matchingBytes[416]),
.io_matchingBytes_417(matchingBytes[417]),
.io_matchingBytes_418(matchingBytes[418]),
.io_matchingBytes_419(matchingBytes[419]),
.io_matchingBytes_420(matchingBytes[420]),
.io_matchingBytes_421(matchingBytes[421]),
.io_matchingBytes_422(matchingBytes[422]),
.io_matchingBytes_423(matchingBytes[423]),
.io_matchingBytes_424(matchingBytes[424]),
.io_matchingBytes_425(matchingBytes[425]),
.io_matchingBytes_426(matchingBytes[426]),
.io_matchingBytes_427(matchingBytes[427]),
.io_matchingBytes_428(matchingBytes[428]),
.io_matchingBytes_429(matchingBytes[429]),
.io_matchingBytes_430(matchingBytes[430]),
.io_matchingBytes_431(matchingBytes[431]),
.io_matchingBytes_432(matchingBytes[432]),
.io_matchingBytes_433(matchingBytes[433]),
.io_matchingBytes_434(matchingBytes[434]),
.io_matchingBytes_435(matchingBytes[435]),
.io_matchingBytes_436(matchingBytes[436]),
.io_matchingBytes_437(matchingBytes[437]),
.io_matchingBytes_438(matchingBytes[438]),
.io_matchingBytes_439(matchingBytes[439]),
.io_matchingBytes_440(matchingBytes[440]),
.io_matchingBytes_441(matchingBytes[441]),
.io_matchingBytes_442(matchingBytes[442]),
.io_matchingBytes_443(matchingBytes[443]),
.io_matchingBytes_444(matchingBytes[444]),
.io_matchingBytes_445(matchingBytes[445]),
.io_matchingBytes_446(matchingBytes[446]),
.io_matchingBytes_447(matchingBytes[447]),
.io_matchingBytes_448(matchingBytes[448]),
.io_matchingBytes_449(matchingBytes[449]),
.io_matchingBytes_450(matchingBytes[450]),
.io_matchingBytes_451(matchingBytes[451]),
.io_matchingBytes_452(matchingBytes[452]),
.io_matchingBytes_453(matchingBytes[453]),
.io_matchingBytes_454(matchingBytes[454]),
.io_matchingBytes_455(matchingBytes[455]),
.io_matchingBytes_456(matchingBytes[456]),
.io_matchingBytes_457(matchingBytes[457]),
.io_matchingBytes_458(matchingBytes[458]),
.io_matchingBytes_459(matchingBytes[459]),
.io_matchingBytes_460(matchingBytes[460]),
.io_matchingBytes_461(matchingBytes[461]),
.io_matchingBytes_462(matchingBytes[462]),
.io_matchingBytes_463(matchingBytes[463]),
.io_matchingBytes_464(matchingBytes[464]),
.io_matchingBytes_465(matchingBytes[465]),
.io_matchingBytes_466(matchingBytes[466]),
.io_matchingBytes_467(matchingBytes[467]),
.io_matchingBytes_468(matchingBytes[468]),
.io_matchingBytes_469(matchingBytes[469]),
.io_matchingBytes_470(matchingBytes[470]),
.io_matchingBytes_471(matchingBytes[471]),
.io_matchingBytes_472(matchingBytes[472]),
.io_matchingBytes_473(matchingBytes[473]),
.io_matchingBytes_474(matchingBytes[474]),
.io_matchingBytes_475(matchingBytes[475]),
.io_matchingBytes_476(matchingBytes[476]),
.io_matchingBytes_477(matchingBytes[477]),
.io_matchingBytes_478(matchingBytes[478]),
.io_matchingBytes_479(matchingBytes[479]),
.io_matchingBytes_480(matchingBytes[480]),
.io_matchingBytes_481(matchingBytes[481]),
.io_matchingBytes_482(matchingBytes[482]),
.io_matchingBytes_483(matchingBytes[483]),
.io_matchingBytes_484(matchingBytes[484]),
.io_matchingBytes_485(matchingBytes[485]),
.io_matchingBytes_486(matchingBytes[486]),
.io_matchingBytes_487(matchingBytes[487]),
.io_matchingBytes_488(matchingBytes[488]),
.io_matchingBytes_489(matchingBytes[489]),
.io_matchingBytes_490(matchingBytes[490]),
.io_matchingBytes_491(matchingBytes[491]),
.io_matchingBytes_492(matchingBytes[492]),
.io_matchingBytes_493(matchingBytes[493]),
.io_matchingBytes_494(matchingBytes[494]),
.io_matchingBytes_495(matchingBytes[495]),
.io_matchingBytes_496(matchingBytes[496]),
.io_matchingBytes_497(matchingBytes[497]),
.io_matchingBytes_498(matchingBytes[498]),
.io_matchingBytes_499(matchingBytes[499]),
.io_matchingBytes_500(matchingBytes[500]),
.io_matchingBytes_501(matchingBytes[501]),
.io_matchingBytes_502(matchingBytes[502]),
.io_matchingBytes_503(matchingBytes[503]),
.io_matchingBytes_504(matchingBytes[504]),
.io_matchingBytes_505(matchingBytes[505]),
.io_matchingBytes_506(matchingBytes[506]),
.io_matchingBytes_507(matchingBytes[507]),
.io_matchingBytes_508(matchingBytes[508]),
.io_matchingBytes_509(matchingBytes[509]),
.io_matchingBytes_510(matchingBytes[510]),
.io_matchingBytes_511(matchingBytes[511]),
.io_matchingBytes_512(matchingBytes[512]),
.io_matchingBytes_513(matchingBytes[513]),
.io_matchingBytes_514(matchingBytes[514]),
.io_matchingBytes_515(matchingBytes[515]),
.io_matchingBytes_516(matchingBytes[516]),
.io_matchingBytes_517(matchingBytes[517]),
.io_matchingBytes_518(matchingBytes[518]),
.io_matchingBytes_519(matchingBytes[519]),
.io_matchingBytes_520(matchingBytes[520]),
.io_matchingBytes_521(matchingBytes[521]),
.io_matchingBytes_522(matchingBytes[522]),
.io_matchingBytes_523(matchingBytes[523]),
.io_matchingBytes_524(matchingBytes[524]),
.io_matchingBytes_525(matchingBytes[525]),
.io_matchingBytes_526(matchingBytes[526]),
.io_matchingBytes_527(matchingBytes[527]),
.io_matchingBytes_528(matchingBytes[528]),
.io_matchingBytes_529(matchingBytes[529]),
.io_matchingBytes_530(matchingBytes[530]),
.io_matchingBytes_531(matchingBytes[531]),
.io_matchingBytes_532(matchingBytes[532]),
.io_matchingBytes_533(matchingBytes[533]),
.io_matchingBytes_534(matchingBytes[534]),
.io_matchingBytes_535(matchingBytes[535]),
.io_matchingBytes_536(matchingBytes[536]),
.io_matchingBytes_537(matchingBytes[537]),
.io_matchingBytes_538(matchingBytes[538]),
.io_matchingBytes_539(matchingBytes[539]),
.io_matchingBytes_540(matchingBytes[540]),
.io_matchingBytes_541(matchingBytes[541]),
.io_matchingBytes_542(matchingBytes[542]),
.io_matchingBytes_543(matchingBytes[543]),
.io_matchingBytes_544(matchingBytes[544]),
.io_matchingBytes_545(matchingBytes[545]),
.io_matchingBytes_546(matchingBytes[546]),
.io_matchingBytes_547(matchingBytes[547]),
.io_matchingBytes_548(matchingBytes[548]),
.io_matchingBytes_549(matchingBytes[549]),
.io_matchingBytes_550(matchingBytes[550]),
.io_matchingBytes_551(matchingBytes[551]),
.io_matchingBytes_552(matchingBytes[552]),
.io_matchingBytes_553(matchingBytes[553]),
.io_matchingBytes_554(matchingBytes[554]),
.io_matchingBytes_555(matchingBytes[555]),
.io_matchingBytes_556(matchingBytes[556]),
.io_matchingBytes_557(matchingBytes[557]),
.io_matchingBytes_558(matchingBytes[558]),
.io_matchingBytes_559(matchingBytes[559]),
.io_matchingBytes_560(matchingBytes[560]),
.io_matchingBytes_561(matchingBytes[561]),
.io_matchingBytes_562(matchingBytes[562]),
.io_matchingBytes_563(matchingBytes[563]),
.io_matchingBytes_564(matchingBytes[564]),
.io_matchingBytes_565(matchingBytes[565]),
.io_matchingBytes_566(matchingBytes[566]),
.io_matchingBytes_567(matchingBytes[567]),
.io_matchingBytes_568(matchingBytes[568]),
.io_matchingBytes_569(matchingBytes[569]),
.io_matchingBytes_570(matchingBytes[570]),
.io_matchingBytes_571(matchingBytes[571]),
.io_matchingBytes_572(matchingBytes[572]),
.io_matchingBytes_573(matchingBytes[573]),
.io_matchingBytes_574(matchingBytes[574]),
.io_matchingBytes_575(matchingBytes[575]),
.io_matchingBytes_576(matchingBytes[576]),
.io_matchingBytes_577(matchingBytes[577]),
.io_matchingBytes_578(matchingBytes[578]),
.io_matchingBytes_579(matchingBytes[579]),
.io_matchingBytes_580(matchingBytes[580]),
.io_matchingBytes_581(matchingBytes[581]),
.io_matchingBytes_582(matchingBytes[582]),
.io_matchingBytes_583(matchingBytes[583]),
.io_matchingBytes_584(matchingBytes[584]),
.io_matchingBytes_585(matchingBytes[585]),
.io_matchingBytes_586(matchingBytes[586]),
.io_matchingBytes_587(matchingBytes[587]),
.io_matchingBytes_588(matchingBytes[588]),
.io_matchingBytes_589(matchingBytes[589]),
.io_matchingBytes_590(matchingBytes[590]),
.io_matchingBytes_591(matchingBytes[591]),
.io_matchingBytes_592(matchingBytes[592]),
.io_matchingBytes_593(matchingBytes[593]),
.io_matchingBytes_594(matchingBytes[594]),
.io_matchingBytes_595(matchingBytes[595]),
.io_matchingBytes_596(matchingBytes[596]),
.io_matchingBytes_597(matchingBytes[597]),
.io_matchingBytes_598(matchingBytes[598]),
.io_matchingBytes_599(matchingBytes[599]),
.io_matchingBytes_600(matchingBytes[600]),
.io_matchingBytes_601(matchingBytes[601]),
.io_matchingBytes_602(matchingBytes[602]),
.io_matchingBytes_603(matchingBytes[603]),
.io_matchingBytes_604(matchingBytes[604]),
.io_matchingBytes_605(matchingBytes[605]),
.io_matchingBytes_606(matchingBytes[606]),
.io_matchingBytes_607(matchingBytes[607]),
.io_matchingBytes_608(matchingBytes[608]),
.io_matchingBytes_609(matchingBytes[609]),
.io_matchingBytes_610(matchingBytes[610]),
.io_matchingBytes_611(matchingBytes[611]),
.io_matchingBytes_612(matchingBytes[612]),
.io_matchingBytes_613(matchingBytes[613]),
.io_matchingBytes_614(matchingBytes[614]),
.io_matchingBytes_615(matchingBytes[615]),
.io_matchingBytes_616(matchingBytes[616]),
.io_matchingBytes_617(matchingBytes[617]),
.io_matchingBytes_618(matchingBytes[618]),
.io_matchingBytes_619(matchingBytes[619]),
.io_matchingBytes_620(matchingBytes[620]),
.io_matchingBytes_621(matchingBytes[621]),
.io_matchingBytes_622(matchingBytes[622]),
.io_matchingBytes_623(matchingBytes[623]),
.io_matchingBytes_624(matchingBytes[624]),
.io_matchingBytes_625(matchingBytes[625]),
.io_matchingBytes_626(matchingBytes[626]),
.io_matchingBytes_627(matchingBytes[627]),
.io_matchingBytes_628(matchingBytes[628]),
.io_matchingBytes_629(matchingBytes[629]),
.io_matchingBytes_630(matchingBytes[630]),
.io_matchingBytes_631(matchingBytes[631]),
.io_matchingBytes_632(matchingBytes[632]),
.io_matchingBytes_633(matchingBytes[633]),
.io_matchingBytes_634(matchingBytes[634]),
.io_matchingBytes_635(matchingBytes[635]),
.io_matchingBytes_636(matchingBytes[636]),
.io_matchingBytes_637(matchingBytes[637]),
.io_matchingBytes_638(matchingBytes[638]),
.io_matchingBytes_639(matchingBytes[639]),
.io_matchingBytes_640(matchingBytes[640]),
.io_matchingBytes_641(matchingBytes[641]),
.io_matchingBytes_642(matchingBytes[642]),
.io_matchingBytes_643(matchingBytes[643]),
.io_matchingBytes_644(matchingBytes[644]),
.io_matchingBytes_645(matchingBytes[645]),
.io_matchingBytes_646(matchingBytes[646]),
.io_matchingBytes_647(matchingBytes[647]),
.io_matchingBytes_648(matchingBytes[648]),
.io_matchingBytes_649(matchingBytes[649]),
.io_matchingBytes_650(matchingBytes[650]),
.io_matchingBytes_651(matchingBytes[651]),
.io_matchingBytes_652(matchingBytes[652]),
.io_matchingBytes_653(matchingBytes[653]),
.io_matchingBytes_654(matchingBytes[654]),
.io_matchingBytes_655(matchingBytes[655]),
.io_matchingBytes_656(matchingBytes[656]),
.io_matchingBytes_657(matchingBytes[657]),
.io_matchingBytes_658(matchingBytes[658]),
.io_matchingBytes_659(matchingBytes[659]),
.io_matchingBytes_660(matchingBytes[660]),
.io_matchingBytes_661(matchingBytes[661]),
.io_matchingBytes_662(matchingBytes[662]),
.io_matchingBytes_663(matchingBytes[663]),
.io_matchingBytes_664(matchingBytes[664]),
.io_matchingBytes_665(matchingBytes[665]),
.io_matchingBytes_666(matchingBytes[666]),
.io_matchingBytes_667(matchingBytes[667]),
.io_matchingBytes_668(matchingBytes[668]),
.io_matchingBytes_669(matchingBytes[669]),
.io_matchingBytes_670(matchingBytes[670]),
.io_matchingBytes_671(matchingBytes[671]),
.io_matchingBytes_672(matchingBytes[672]),
.io_matchingBytes_673(matchingBytes[673]),
.io_matchingBytes_674(matchingBytes[674]),
.io_matchingBytes_675(matchingBytes[675]),
.io_matchingBytes_676(matchingBytes[676]),
.io_matchingBytes_677(matchingBytes[677]),
.io_matchingBytes_678(matchingBytes[678]),
.io_matchingBytes_679(matchingBytes[679]),
.io_matchingBytes_680(matchingBytes[680]),
.io_matchingBytes_681(matchingBytes[681]),
.io_matchingBytes_682(matchingBytes[682]),
.io_matchingBytes_683(matchingBytes[683]),
.io_matchingBytes_684(matchingBytes[684]),
.io_matchingBytes_685(matchingBytes[685]),
.io_matchingBytes_686(matchingBytes[686]),
.io_matchingBytes_687(matchingBytes[687]),
.io_matchingBytes_688(matchingBytes[688]),
.io_matchingBytes_689(matchingBytes[689]),
.io_matchingBytes_690(matchingBytes[690]),
.io_matchingBytes_691(matchingBytes[691]),
.io_matchingBytes_692(matchingBytes[692]),
.io_matchingBytes_693(matchingBytes[693]),
.io_matchingBytes_694(matchingBytes[694]),
.io_matchingBytes_695(matchingBytes[695]),
.io_matchingBytes_696(matchingBytes[696]),
.io_matchingBytes_697(matchingBytes[697]),
.io_matchingBytes_698(matchingBytes[698]),
.io_matchingBytes_699(matchingBytes[699]),
.io_matchingBytes_700(matchingBytes[700]),
.io_matchingBytes_701(matchingBytes[701]),
.io_matchingBytes_702(matchingBytes[702]),
.io_matchingBytes_703(matchingBytes[703]),
.io_matchingBytes_704(matchingBytes[704]),
.io_matchingBytes_705(matchingBytes[705]),
.io_matchingBytes_706(matchingBytes[706]),
.io_matchingBytes_707(matchingBytes[707]),
.io_matchingBytes_708(matchingBytes[708]),
.io_matchingBytes_709(matchingBytes[709]),
.io_matchingBytes_710(matchingBytes[710]),
.io_matchingBytes_711(matchingBytes[711]),
.io_matchingBytes_712(matchingBytes[712]),
.io_matchingBytes_713(matchingBytes[713]),
.io_matchingBytes_714(matchingBytes[714]),
.io_matchingBytes_715(matchingBytes[715]),
.io_matchingBytes_716(matchingBytes[716]),
.io_matchingBytes_717(matchingBytes[717]),
.io_matchingBytes_718(matchingBytes[718]),
.io_matchingBytes_719(matchingBytes[719]),
.io_matchingBytes_720(matchingBytes[720]),
.io_matchingBytes_721(matchingBytes[721]),
.io_matchingBytes_722(matchingBytes[722]),
.io_matchingBytes_723(matchingBytes[723]),
.io_matchingBytes_724(matchingBytes[724]),
.io_matchingBytes_725(matchingBytes[725]),
.io_matchingBytes_726(matchingBytes[726]),
.io_matchingBytes_727(matchingBytes[727]),
.io_matchingBytes_728(matchingBytes[728]),
.io_matchingBytes_729(matchingBytes[729]),
.io_matchingBytes_730(matchingBytes[730]),
.io_matchingBytes_731(matchingBytes[731]),
.io_matchingBytes_732(matchingBytes[732]),
.io_matchingBytes_733(matchingBytes[733]),
.io_matchingBytes_734(matchingBytes[734]),
.io_matchingBytes_735(matchingBytes[735]),
.io_matchingBytes_736(matchingBytes[736]),
.io_matchingBytes_737(matchingBytes[737]),
.io_matchingBytes_738(matchingBytes[738]),
.io_matchingBytes_739(matchingBytes[739]),
.io_matchingBytes_740(matchingBytes[740]),
.io_matchingBytes_741(matchingBytes[741]),
.io_matchingBytes_742(matchingBytes[742]),
.io_matchingBytes_743(matchingBytes[743]),
.io_matchingBytes_744(matchingBytes[744]),
.io_matchingBytes_745(matchingBytes[745]),
.io_matchingBytes_746(matchingBytes[746]),
.io_matchingBytes_747(matchingBytes[747]),
.io_matchingBytes_748(matchingBytes[748]),
.io_matchingBytes_749(matchingBytes[749]),
.io_matchingBytes_750(matchingBytes[750]),
.io_matchingBytes_751(matchingBytes[751]),
.io_matchingBytes_752(matchingBytes[752]),
.io_matchingBytes_753(matchingBytes[753]),
.io_matchingBytes_754(matchingBytes[754]),
.io_matchingBytes_755(matchingBytes[755]),
.io_matchingBytes_756(matchingBytes[756]),
.io_matchingBytes_757(matchingBytes[757]),
.io_matchingBytes_758(matchingBytes[758]),
.io_matchingBytes_759(matchingBytes[759]),
.io_matchingBytes_760(matchingBytes[760]),
.io_matchingBytes_761(matchingBytes[761]),
.io_matchingBytes_762(matchingBytes[762]),
.io_matchingBytes_763(matchingBytes[763]),
.io_matchingBytes_764(matchingBytes[764]),
.io_matchingBytes_765(matchingBytes[765]),
.io_matchingBytes_766(matchingBytes[766]),
.io_matchingBytes_767(matchingBytes[767]),
.io_matchingBytes_768(matchingBytes[768]),
.io_matchingBytes_769(matchingBytes[769]),
.io_matchingBytes_770(matchingBytes[770]),
.io_matchingBytes_771(matchingBytes[771]),
.io_matchingBytes_772(matchingBytes[772]),
.io_matchingBytes_773(matchingBytes[773]),
.io_matchingBytes_774(matchingBytes[774]),
.io_matchingBytes_775(matchingBytes[775]),
.io_matchingBytes_776(matchingBytes[776]),
.io_matchingBytes_777(matchingBytes[777]),
.io_matchingBytes_778(matchingBytes[778]),
.io_matchingBytes_779(matchingBytes[779]),
.io_matchingBytes_780(matchingBytes[780]),
.io_matchingBytes_781(matchingBytes[781]),
.io_matchingBytes_782(matchingBytes[782]),
.io_matchingBytes_783(matchingBytes[783]),
.io_matchingBytes_784(matchingBytes[784]),
.io_matchingBytes_785(matchingBytes[785]),
.io_matchingBytes_786(matchingBytes[786]),
.io_matchingBytes_787(matchingBytes[787]),
.io_matchingBytes_788(matchingBytes[788]),
.io_matchingBytes_789(matchingBytes[789]),
.io_matchingBytes_790(matchingBytes[790]),
.io_matchingBytes_791(matchingBytes[791]),
.io_matchingBytes_792(matchingBytes[792]),
.io_matchingBytes_793(matchingBytes[793]),
.io_matchingBytes_794(matchingBytes[794]),
.io_matchingBytes_795(matchingBytes[795]),
.io_matchingBytes_796(matchingBytes[796]),
.io_matchingBytes_797(matchingBytes[797]),
.io_matchingBytes_798(matchingBytes[798]),
.io_matchingBytes_799(matchingBytes[799]),
.io_matchingBytes_800(matchingBytes[800]),
.io_matchingBytes_801(matchingBytes[801]),
.io_matchingBytes_802(matchingBytes[802]),
.io_matchingBytes_803(matchingBytes[803]),
.io_matchingBytes_804(matchingBytes[804]),
.io_matchingBytes_805(matchingBytes[805]),
.io_matchingBytes_806(matchingBytes[806]),
.io_matchingBytes_807(matchingBytes[807]),
.io_matchingBytes_808(matchingBytes[808]),
.io_matchingBytes_809(matchingBytes[809]),
.io_matchingBytes_810(matchingBytes[810]),
.io_matchingBytes_811(matchingBytes[811]),
.io_matchingBytes_812(matchingBytes[812]),
.io_matchingBytes_813(matchingBytes[813]),
.io_matchingBytes_814(matchingBytes[814]),
.io_matchingBytes_815(matchingBytes[815]),
.io_matchingBytes_816(matchingBytes[816]),
.io_matchingBytes_817(matchingBytes[817]),
.io_matchingBytes_818(matchingBytes[818]),
.io_matchingBytes_819(matchingBytes[819]),
.io_matchingBytes_820(matchingBytes[820]),
.io_matchingBytes_821(matchingBytes[821]),
.io_matchingBytes_822(matchingBytes[822]),
.io_matchingBytes_823(matchingBytes[823]),
.io_matchingBytes_824(matchingBytes[824]),
.io_matchingBytes_825(matchingBytes[825]),
.io_matchingBytes_826(matchingBytes[826]),
.io_matchingBytes_827(matchingBytes[827]),
.io_matchingBytes_828(matchingBytes[828]),
.io_matchingBytes_829(matchingBytes[829]),
.io_matchingBytes_830(matchingBytes[830]),
.io_matchingBytes_831(matchingBytes[831]),
.io_matchingBytes_832(matchingBytes[832]),
.io_matchingBytes_833(matchingBytes[833]),
.io_matchingBytes_834(matchingBytes[834]),
.io_matchingBytes_835(matchingBytes[835]),
.io_matchingBytes_836(matchingBytes[836]),
.io_matchingBytes_837(matchingBytes[837]),
.io_matchingBytes_838(matchingBytes[838]),
.io_matchingBytes_839(matchingBytes[839]),
.io_matchingBytes_840(matchingBytes[840]),
.io_matchingBytes_841(matchingBytes[841]),
.io_matchingBytes_842(matchingBytes[842]),
.io_matchingBytes_843(matchingBytes[843]),
.io_matchingBytes_844(matchingBytes[844]),
.io_matchingBytes_845(matchingBytes[845]),
.io_matchingBytes_846(matchingBytes[846]),
.io_matchingBytes_847(matchingBytes[847]),
.io_matchingBytes_848(matchingBytes[848]),
.io_matchingBytes_849(matchingBytes[849]),
.io_matchingBytes_850(matchingBytes[850]),
.io_matchingBytes_851(matchingBytes[851]),
.io_matchingBytes_852(matchingBytes[852]),
.io_matchingBytes_853(matchingBytes[853]),
.io_matchingBytes_854(matchingBytes[854]),
.io_matchingBytes_855(matchingBytes[855]),
.io_matchingBytes_856(matchingBytes[856]),
.io_matchingBytes_857(matchingBytes[857]),
.io_matchingBytes_858(matchingBytes[858]),
.io_matchingBytes_859(matchingBytes[859]),
.io_matchingBytes_860(matchingBytes[860]),
.io_matchingBytes_861(matchingBytes[861]),
.io_matchingBytes_862(matchingBytes[862]),
.io_matchingBytes_863(matchingBytes[863]),
.io_matchingBytes_864(matchingBytes[864]),
.io_matchingBytes_865(matchingBytes[865]),
.io_matchingBytes_866(matchingBytes[866]),
.io_matchingBytes_867(matchingBytes[867]),
.io_matchingBytes_868(matchingBytes[868]),
.io_matchingBytes_869(matchingBytes[869]),
.io_matchingBytes_870(matchingBytes[870]),
.io_matchingBytes_871(matchingBytes[871]),
.io_matchingBytes_872(matchingBytes[872]),
.io_matchingBytes_873(matchingBytes[873]),
.io_matchingBytes_874(matchingBytes[874]),
.io_matchingBytes_875(matchingBytes[875]),
.io_matchingBytes_876(matchingBytes[876]),
.io_matchingBytes_877(matchingBytes[877]),
.io_matchingBytes_878(matchingBytes[878]),
.io_matchingBytes_879(matchingBytes[879]),
.io_matchingBytes_880(matchingBytes[880]),
.io_matchingBytes_881(matchingBytes[881]),
.io_matchingBytes_882(matchingBytes[882]),
.io_matchingBytes_883(matchingBytes[883]),
.io_matchingBytes_884(matchingBytes[884]),
.io_matchingBytes_885(matchingBytes[885]),
.io_matchingBytes_886(matchingBytes[886]),
.io_matchingBytes_887(matchingBytes[887]),
.io_matchingBytes_888(matchingBytes[888]),
.io_matchingBytes_889(matchingBytes[889]),
.io_matchingBytes_890(matchingBytes[890]),
.io_matchingBytes_891(matchingBytes[891]),
.io_matchingBytes_892(matchingBytes[892]),
.io_matchingBytes_893(matchingBytes[893]),
.io_matchingBytes_894(matchingBytes[894]),
.io_matchingBytes_895(matchingBytes[895]),
.io_matchingBytes_896(matchingBytes[896]),
.io_matchingBytes_897(matchingBytes[897]),
.io_matchingBytes_898(matchingBytes[898]),
.io_matchingBytes_899(matchingBytes[899]),
.io_matchingBytes_900(matchingBytes[900]),
.io_matchingBytes_901(matchingBytes[901]),
.io_matchingBytes_902(matchingBytes[902]),
.io_matchingBytes_903(matchingBytes[903]),
.io_matchingBytes_904(matchingBytes[904]),
.io_matchingBytes_905(matchingBytes[905]),
.io_matchingBytes_906(matchingBytes[906]),
.io_matchingBytes_907(matchingBytes[907]),
.io_matchingBytes_908(matchingBytes[908]),
.io_matchingBytes_909(matchingBytes[909]),
.io_matchingBytes_910(matchingBytes[910]),
.io_matchingBytes_911(matchingBytes[911]),
.io_matchingBytes_912(matchingBytes[912]),
.io_matchingBytes_913(matchingBytes[913]),
.io_matchingBytes_914(matchingBytes[914]),
.io_matchingBytes_915(matchingBytes[915]),
.io_matchingBytes_916(matchingBytes[916]),
.io_matchingBytes_917(matchingBytes[917]),
.io_matchingBytes_918(matchingBytes[918]),
.io_matchingBytes_919(matchingBytes[919]),
.io_matchingBytes_920(matchingBytes[920]),
.io_matchingBytes_921(matchingBytes[921]),
.io_matchingBytes_922(matchingBytes[922]),
.io_matchingBytes_923(matchingBytes[923]),
.io_matchingBytes_924(matchingBytes[924]),
.io_matchingBytes_925(matchingBytes[925]),
.io_matchingBytes_926(matchingBytes[926]),
.io_matchingBytes_927(matchingBytes[927]),
.io_matchingBytes_928(matchingBytes[928]),
.io_matchingBytes_929(matchingBytes[929]),
.io_matchingBytes_930(matchingBytes[930]),
.io_matchingBytes_931(matchingBytes[931]),
.io_matchingBytes_932(matchingBytes[932]),
.io_matchingBytes_933(matchingBytes[933]),
.io_matchingBytes_934(matchingBytes[934]),
.io_matchingBytes_935(matchingBytes[935]),
.io_matchingBytes_936(matchingBytes[936]),
.io_matchingBytes_937(matchingBytes[937]),
.io_matchingBytes_938(matchingBytes[938]),
.io_matchingBytes_939(matchingBytes[939]),
.io_matchingBytes_940(matchingBytes[940]),
.io_matchingBytes_941(matchingBytes[941]),
.io_matchingBytes_942(matchingBytes[942]),
.io_matchingBytes_943(matchingBytes[943]),
.io_matchingBytes_944(matchingBytes[944]),
.io_matchingBytes_945(matchingBytes[945]),
.io_matchingBytes_946(matchingBytes[946]),
.io_matchingBytes_947(matchingBytes[947]),
.io_matchingBytes_948(matchingBytes[948]),
.io_matchingBytes_949(matchingBytes[949]),
.io_matchingBytes_950(matchingBytes[950]),
.io_matchingBytes_951(matchingBytes[951]),
.io_matchingBytes_952(matchingBytes[952]),
.io_matchingBytes_953(matchingBytes[953]),
.io_matchingBytes_954(matchingBytes[954]),
.io_matchingBytes_955(matchingBytes[955]),
.io_matchingBytes_956(matchingBytes[956]),
.io_matchingBytes_957(matchingBytes[957]),
.io_matchingBytes_958(matchingBytes[958]),
.io_matchingBytes_959(matchingBytes[959]),
.io_matchingBytes_960(matchingBytes[960]),
.io_matchingBytes_961(matchingBytes[961]),
.io_matchingBytes_962(matchingBytes[962]),
.io_matchingBytes_963(matchingBytes[963]),
.io_matchingBytes_964(matchingBytes[964]),
.io_matchingBytes_965(matchingBytes[965]),
.io_matchingBytes_966(matchingBytes[966]),
.io_matchingBytes_967(matchingBytes[967]),
.io_matchingBytes_968(matchingBytes[968]),
.io_matchingBytes_969(matchingBytes[969]),
.io_matchingBytes_970(matchingBytes[970]),
.io_matchingBytes_971(matchingBytes[971]),
.io_matchingBytes_972(matchingBytes[972]),
.io_matchingBytes_973(matchingBytes[973]),
.io_matchingBytes_974(matchingBytes[974]),
.io_matchingBytes_975(matchingBytes[975]),
.io_matchingBytes_976(matchingBytes[976]),
.io_matchingBytes_977(matchingBytes[977]),
.io_matchingBytes_978(matchingBytes[978]),
.io_matchingBytes_979(matchingBytes[979]),
.io_matchingBytes_980(matchingBytes[980]),
.io_matchingBytes_981(matchingBytes[981]),
.io_matchingBytes_982(matchingBytes[982]),
.io_matchingBytes_983(matchingBytes[983]),
.io_matchingBytes_984(matchingBytes[984]),
.io_matchingBytes_985(matchingBytes[985]),
.io_matchingBytes_986(matchingBytes[986]),
.io_matchingBytes_987(matchingBytes[987]),
.io_matchingBytes_988(matchingBytes[988]),
.io_matchingBytes_989(matchingBytes[989]),
.io_matchingBytes_990(matchingBytes[990]),
.io_matchingBytes_991(matchingBytes[991]),
.io_matchingBytes_992(matchingBytes[992]),
.io_matchingBytes_993(matchingBytes[993]),
.io_matchingBytes_994(matchingBytes[994]),
.io_matchingBytes_995(matchingBytes[995]),
.io_matchingBytes_996(matchingBytes[996]),
.io_matchingBytes_997(matchingBytes[997]),
.io_matchingBytes_998(matchingBytes[998]),
.io_matchingBytes_999(matchingBytes[999]),
.io_matchingBytes_1000(matchingBytes[1000]),
.io_matchingBytes_1001(matchingBytes[1001]),
.io_matchingBytes_1002(matchingBytes[1002]),
.io_matchingBytes_1003(matchingBytes[1003]),
.io_matchingBytes_1004(matchingBytes[1004]),
.io_matchingBytes_1005(matchingBytes[1005]),
.io_matchingBytes_1006(matchingBytes[1006]),
.io_matchingBytes_1007(matchingBytes[1007]),
.io_matchingBytes_1008(matchingBytes[1008]),
.io_matchingBytes_1009(matchingBytes[1009]),
.io_matchingBytes_1010(matchingBytes[1010]),
.io_matchingBytes_1011(matchingBytes[1011]),
.io_matchingBytes_1012(matchingBytes[1012]),
.io_matchingBytes_1013(matchingBytes[1013]),
.io_matchingBytes_1014(matchingBytes[1014]),
.io_matchingBytes_1015(matchingBytes[1015]),
.io_matchingBytes_1016(matchingBytes[1016]),
.io_matchingBytes_1017(matchingBytes[1017]),
.io_matchingBytes_1018(matchingBytes[1018]),
.io_matchingBytes_1019(matchingBytes[1019]),
.io_matchingBytes_1020(matchingBytes[1020]),
.io_matchingBytes_1021(matchingBytes[1021]),
.io_matchingBytes_1022(matchingBytes[1022]),
.io_matchingBytes_1023(matchingBytes[1023]),
.io_matchingBytes_1024(matchingBytes[1024]),
.io_matchingBytes_1025(matchingBytes[1025]),
.io_matchingBytes_1026(matchingBytes[1026]),
.io_matchingBytes_1027(matchingBytes[1027]),
.io_matchingBytes_1028(matchingBytes[1028]),
.io_matchingBytes_1029(matchingBytes[1029]),
.io_matchingBytes_1030(matchingBytes[1030]),
.io_matchingBytes_1031(matchingBytes[1031]),
.io_matchingBytes_1032(matchingBytes[1032]),
.io_matchingBytes_1033(matchingBytes[1033]),
.io_matchingBytes_1034(matchingBytes[1034]),
.io_matchingBytes_1035(matchingBytes[1035]),
.io_matchingBytes_1036(matchingBytes[1036]),
.io_matchingBytes_1037(matchingBytes[1037]),
.io_matchingBytes_1038(matchingBytes[1038]),
.io_matchingBytes_1039(matchingBytes[1039]),
.io_matchingBytes_1040(matchingBytes[1040]),
.io_matchingBytes_1041(matchingBytes[1041]),
.io_matchingBytes_1042(matchingBytes[1042]),
.io_matchingBytes_1043(matchingBytes[1043]),
.io_matchingBytes_1044(matchingBytes[1044]),
.io_matchingBytes_1045(matchingBytes[1045]),
.io_matchingBytes_1046(matchingBytes[1046]),
.io_matchingBytes_1047(matchingBytes[1047]),
.io_matchingBytes_1048(matchingBytes[1048]),
.io_matchingBytes_1049(matchingBytes[1049]),
.io_matchingBytes_1050(matchingBytes[1050]),
.io_matchingBytes_1051(matchingBytes[1051]),
.io_matchingBytes_1052(matchingBytes[1052]),
.io_matchingBytes_1053(matchingBytes[1053]),
.io_matchingBytes_1054(matchingBytes[1054]),
.io_matchingBytes_1055(matchingBytes[1055]),
.io_matchingBytes_1056(matchingBytes[1056]),
.io_matchingBytes_1057(matchingBytes[1057]),
.io_matchingBytes_1058(matchingBytes[1058]),
.io_matchingBytes_1059(matchingBytes[1059]),
.io_matchingBytes_1060(matchingBytes[1060]),
.io_matchingBytes_1061(matchingBytes[1061]),
.io_matchingBytes_1062(matchingBytes[1062]),
.io_matchingBytes_1063(matchingBytes[1063]),
.io_matchingBytes_1064(matchingBytes[1064]),
.io_matchingBytes_1065(matchingBytes[1065]),
.io_matchingBytes_1066(matchingBytes[1066]),
.io_matchingBytes_1067(matchingBytes[1067]),
.io_matchingBytes_1068(matchingBytes[1068]),
.io_matchingBytes_1069(matchingBytes[1069]),
.io_matchingBytes_1070(matchingBytes[1070]),
.io_matchingBytes_1071(matchingBytes[1071]),
.io_matchingBytes_1072(matchingBytes[1072]),
.io_matchingBytes_1073(matchingBytes[1073]),
.io_matchingBytes_1074(matchingBytes[1074]),
.io_matchingBytes_1075(matchingBytes[1075]),
.io_matchingBytes_1076(matchingBytes[1076]),
.io_matchingBytes_1077(matchingBytes[1077]),
.io_matchingBytes_1078(matchingBytes[1078]),
.io_matchingBytes_1079(matchingBytes[1079]),
.io_matchingBytes_1080(matchingBytes[1080]),
.io_matchingBytes_1081(matchingBytes[1081]),
.io_matchingBytes_1082(matchingBytes[1082]),
.io_matchingBytes_1083(matchingBytes[1083]),
.io_matchingBytes_1084(matchingBytes[1084]),
.io_matchingBytes_1085(matchingBytes[1085]),
.io_matchingBytes_1086(matchingBytes[1086]),
.io_matchingBytes_1087(matchingBytes[1087]),
.io_matchingBytes_1088(matchingBytes[1088]),
.io_matchingBytes_1089(matchingBytes[1089]),
.io_matchingBytes_1090(matchingBytes[1090]),
.io_matchingBytes_1091(matchingBytes[1091]),
.io_matchingBytes_1092(matchingBytes[1092]),
.io_matchingBytes_1093(matchingBytes[1093]),
.io_matchingBytes_1094(matchingBytes[1094]),
.io_matchingBytes_1095(matchingBytes[1095]),
.io_matchingBytes_1096(matchingBytes[1096]),
.io_matchingBytes_1097(matchingBytes[1097]),
.io_matchingBytes_1098(matchingBytes[1098]),
.io_matchingBytes_1099(matchingBytes[1099]),
.io_matchingBytes_1100(matchingBytes[1100]),
.io_matchingBytes_1101(matchingBytes[1101]),
.io_matchingBytes_1102(matchingBytes[1102]),
.io_matchingBytes_1103(matchingBytes[1103]),
.io_matchingBytes_1104(matchingBytes[1104]),
.io_matchingBytes_1105(matchingBytes[1105]),
.io_matchingBytes_1106(matchingBytes[1106]),
.io_matchingBytes_1107(matchingBytes[1107]),
.io_matchingBytes_1108(matchingBytes[1108]),
.io_matchingBytes_1109(matchingBytes[1109]),
.io_matchingBytes_1110(matchingBytes[1110]),
.io_matchingBytes_1111(matchingBytes[1111]),
.io_matchingBytes_1112(matchingBytes[1112]),
.io_matchingBytes_1113(matchingBytes[1113]),
.io_matchingBytes_1114(matchingBytes[1114]),
.io_matchingBytes_1115(matchingBytes[1115]),
.io_matchingBytes_1116(matchingBytes[1116]),
.io_matchingBytes_1117(matchingBytes[1117]),
.io_matchingBytes_1118(matchingBytes[1118]),
.io_matchingBytes_1119(matchingBytes[1119]),
.io_matchingBytes_1120(matchingBytes[1120]),
.io_matchingBytes_1121(matchingBytes[1121]),
.io_matchingBytes_1122(matchingBytes[1122]),
.io_matchingBytes_1123(matchingBytes[1123]),
.io_matchingBytes_1124(matchingBytes[1124]),
.io_matchingBytes_1125(matchingBytes[1125]),
.io_matchingBytes_1126(matchingBytes[1126]),
.io_matchingBytes_1127(matchingBytes[1127]),
.io_matchingBytes_1128(matchingBytes[1128]),
.io_matchingBytes_1129(matchingBytes[1129]),
.io_matchingBytes_1130(matchingBytes[1130]),
.io_matchingBytes_1131(matchingBytes[1131]),
.io_matchingBytes_1132(matchingBytes[1132]),
.io_matchingBytes_1133(matchingBytes[1133]),
.io_matchingBytes_1134(matchingBytes[1134]),
.io_matchingBytes_1135(matchingBytes[1135]),
.io_matchingBytes_1136(matchingBytes[1136]),
.io_matchingBytes_1137(matchingBytes[1137]),
.io_matchingBytes_1138(matchingBytes[1138]),
.io_matchingBytes_1139(matchingBytes[1139]),
.io_matchingBytes_1140(matchingBytes[1140]),
.io_matchingBytes_1141(matchingBytes[1141]),
.io_matchingBytes_1142(matchingBytes[1142]),
.io_matchingBytes_1143(matchingBytes[1143]),
.io_matchingBytes_1144(matchingBytes[1144]),
.io_matchingBytes_1145(matchingBytes[1145]),
.io_matchingBytes_1146(matchingBytes[1146]),
.io_matchingBytes_1147(matchingBytes[1147]),
.io_matchingBytes_1148(matchingBytes[1148]),
.io_matchingBytes_1149(matchingBytes[1149]),
.io_matchingBytes_1150(matchingBytes[1150]),
.io_matchingBytes_1151(matchingBytes[1151]),
.io_matchingBytes_1152(matchingBytes[1152]),
.io_matchingBytes_1153(matchingBytes[1153]),
.io_matchingBytes_1154(matchingBytes[1154]),
.io_matchingBytes_1155(matchingBytes[1155]),
.io_matchingBytes_1156(matchingBytes[1156]),
.io_matchingBytes_1157(matchingBytes[1157]),
.io_matchingBytes_1158(matchingBytes[1158]),
.io_matchingBytes_1159(matchingBytes[1159]),
.io_matchingBytes_1160(matchingBytes[1160]),
.io_matchingBytes_1161(matchingBytes[1161]),
.io_matchingBytes_1162(matchingBytes[1162]),
.io_matchingBytes_1163(matchingBytes[1163]),
.io_matchingBytes_1164(matchingBytes[1164]),
.io_matchingBytes_1165(matchingBytes[1165]),
.io_matchingBytes_1166(matchingBytes[1166]),
.io_matchingBytes_1167(matchingBytes[1167]),
.io_matchingBytes_1168(matchingBytes[1168]),
.io_matchingBytes_1169(matchingBytes[1169]),
.io_matchingBytes_1170(matchingBytes[1170]),
.io_matchingBytes_1171(matchingBytes[1171]),
.io_matchingBytes_1172(matchingBytes[1172]),
.io_matchingBytes_1173(matchingBytes[1173]),
.io_matchingBytes_1174(matchingBytes[1174]),
.io_matchingBytes_1175(matchingBytes[1175]),
.io_matchingBytes_1176(matchingBytes[1176]),
.io_matchingBytes_1177(matchingBytes[1177]),
.io_matchingBytes_1178(matchingBytes[1178]),
.io_matchingBytes_1179(matchingBytes[1179]),
.io_matchingBytes_1180(matchingBytes[1180]),
.io_matchingBytes_1181(matchingBytes[1181]),
.io_matchingBytes_1182(matchingBytes[1182]),
.io_matchingBytes_1183(matchingBytes[1183]),
.io_matchingBytes_1184(matchingBytes[1184]),
.io_matchingBytes_1185(matchingBytes[1185]),
.io_matchingBytes_1186(matchingBytes[1186]),
.io_matchingBytes_1187(matchingBytes[1187]),
.io_matchingBytes_1188(matchingBytes[1188]),
.io_matchingBytes_1189(matchingBytes[1189]),
.io_matchingBytes_1190(matchingBytes[1190]),
.io_matchingBytes_1191(matchingBytes[1191]),
.io_matchingBytes_1192(matchingBytes[1192]),
.io_matchingBytes_1193(matchingBytes[1193]),
.io_matchingBytes_1194(matchingBytes[1194]),
.io_matchingBytes_1195(matchingBytes[1195]),
.io_matchingBytes_1196(matchingBytes[1196]),
.io_matchingBytes_1197(matchingBytes[1197]),
.io_matchingBytes_1198(matchingBytes[1198]),
.io_matchingBytes_1199(matchingBytes[1199]),
.io_matchingBytes_1200(matchingBytes[1200]),
.io_matchingBytes_1201(matchingBytes[1201]),
.io_matchingBytes_1202(matchingBytes[1202]),
.io_matchingBytes_1203(matchingBytes[1203]),
.io_matchingBytes_1204(matchingBytes[1204]),
.io_matchingBytes_1205(matchingBytes[1205]),
.io_matchingBytes_1206(matchingBytes[1206]),
.io_matchingBytes_1207(matchingBytes[1207]),
.io_matchingBytes_1208(matchingBytes[1208]),
.io_matchingBytes_1209(matchingBytes[1209]),
.io_matchingBytes_1210(matchingBytes[1210]),
.io_matchingBytes_1211(matchingBytes[1211]),
.io_matchingBytes_1212(matchingBytes[1212]),
.io_matchingBytes_1213(matchingBytes[1213]),
.io_matchingBytes_1214(matchingBytes[1214]),
.io_matchingBytes_1215(matchingBytes[1215]),
.io_matchingBytes_1216(matchingBytes[1216]),
.io_matchingBytes_1217(matchingBytes[1217]),
.io_matchingBytes_1218(matchingBytes[1218]),
.io_matchingBytes_1219(matchingBytes[1219]),
.io_matchingBytes_1220(matchingBytes[1220]),
.io_matchingBytes_1221(matchingBytes[1221]),
.io_matchingBytes_1222(matchingBytes[1222]),
.io_matchingBytes_1223(matchingBytes[1223]),
.io_matchingBytes_1224(matchingBytes[1224]),
.io_matchingBytes_1225(matchingBytes[1225]),
.io_matchingBytes_1226(matchingBytes[1226]),
.io_matchingBytes_1227(matchingBytes[1227]),
.io_matchingBytes_1228(matchingBytes[1228]),
.io_matchingBytes_1229(matchingBytes[1229]),
.io_matchingBytes_1230(matchingBytes[1230]),
.io_matchingBytes_1231(matchingBytes[1231]),
.io_matchingBytes_1232(matchingBytes[1232]),
.io_matchingBytes_1233(matchingBytes[1233]),
.io_matchingBytes_1234(matchingBytes[1234]),
.io_matchingBytes_1235(matchingBytes[1235]),
.io_matchingBytes_1236(matchingBytes[1236]),
.io_matchingBytes_1237(matchingBytes[1237]),
.io_matchingBytes_1238(matchingBytes[1238]),
.io_matchingBytes_1239(matchingBytes[1239]),
.io_matchingBytes_1240(matchingBytes[1240]),
.io_matchingBytes_1241(matchingBytes[1241]),
.io_matchingBytes_1242(matchingBytes[1242]),
.io_matchingBytes_1243(matchingBytes[1243]),
.io_matchingBytes_1244(matchingBytes[1244]),
.io_matchingBytes_1245(matchingBytes[1245]),
.io_matchingBytes_1246(matchingBytes[1246]),
.io_matchingBytes_1247(matchingBytes[1247]),
.io_matchingBytes_1248(matchingBytes[1248]),
.io_matchingBytes_1249(matchingBytes[1249]),
.io_matchingBytes_1250(matchingBytes[1250]),
.io_matchingBytes_1251(matchingBytes[1251]),
.io_matchingBytes_1252(matchingBytes[1252]),
.io_matchingBytes_1253(matchingBytes[1253]),
.io_matchingBytes_1254(matchingBytes[1254]),
.io_matchingBytes_1255(matchingBytes[1255]),
.io_matchingBytes_1256(matchingBytes[1256]),
.io_matchingBytes_1257(matchingBytes[1257]),
.io_matchingBytes_1258(matchingBytes[1258]),
.io_matchingBytes_1259(matchingBytes[1259]),
.io_matchingBytes_1260(matchingBytes[1260]),
.io_matchingBytes_1261(matchingBytes[1261]),
.io_matchingBytes_1262(matchingBytes[1262]),
.io_matchingBytes_1263(matchingBytes[1263]),
.io_matchingBytes_1264(matchingBytes[1264]),
.io_matchingBytes_1265(matchingBytes[1265]),
.io_matchingBytes_1266(matchingBytes[1266]),
.io_matchingBytes_1267(matchingBytes[1267]),
.io_matchingBytes_1268(matchingBytes[1268]),
.io_matchingBytes_1269(matchingBytes[1269]),
.io_matchingBytes_1270(matchingBytes[1270]),
.io_matchingBytes_1271(matchingBytes[1271]),
.io_matchingBytes_1272(matchingBytes[1272]),
.io_matchingBytes_1273(matchingBytes[1273]),
.io_matchingBytes_1274(matchingBytes[1274]),
.io_matchingBytes_1275(matchingBytes[1275]),
.io_matchingBytes_1276(matchingBytes[1276]),
.io_matchingBytes_1277(matchingBytes[1277]),
.io_matchingBytes_1278(matchingBytes[1278]),
.io_matchingBytes_1279(matchingBytes[1279]),
.io_matchingBytes_1280(matchingBytes[1280]),
.io_matchingBytes_1281(matchingBytes[1281]),
.io_matchingBytes_1282(matchingBytes[1282]),
.io_matchingBytes_1283(matchingBytes[1283]),
.io_matchingBytes_1284(matchingBytes[1284]),
.io_matchingBytes_1285(matchingBytes[1285]),
.io_matchingBytes_1286(matchingBytes[1286]),
.io_matchingBytes_1287(matchingBytes[1287]),
.io_matchingBytes_1288(matchingBytes[1288]),
.io_matchingBytes_1289(matchingBytes[1289]),
.io_matchingBytes_1290(matchingBytes[1290]),
.io_matchingBytes_1291(matchingBytes[1291]),
.io_matchingBytes_1292(matchingBytes[1292]),
.io_matchingBytes_1293(matchingBytes[1293]),
.io_matchingBytes_1294(matchingBytes[1294]),
.io_matchingBytes_1295(matchingBytes[1295]),
.io_matchingBytes_1296(matchingBytes[1296]),
.io_matchingBytes_1297(matchingBytes[1297]),
.io_matchingBytes_1298(matchingBytes[1298]),
.io_matchingBytes_1299(matchingBytes[1299]),
.io_matchingBytes_1300(matchingBytes[1300]),
.io_matchingBytes_1301(matchingBytes[1301]),
.io_matchingBytes_1302(matchingBytes[1302]),
.io_matchingBytes_1303(matchingBytes[1303]),
.io_matchingBytes_1304(matchingBytes[1304]),
.io_matchingBytes_1305(matchingBytes[1305]),
.io_matchingBytes_1306(matchingBytes[1306]),
.io_matchingBytes_1307(matchingBytes[1307]),
.io_matchingBytes_1308(matchingBytes[1308]),
.io_matchingBytes_1309(matchingBytes[1309]),
.io_matchingBytes_1310(matchingBytes[1310]),
.io_matchingBytes_1311(matchingBytes[1311]),
.io_matchingBytes_1312(matchingBytes[1312]),
.io_matchingBytes_1313(matchingBytes[1313]),
.io_matchingBytes_1314(matchingBytes[1314]),
.io_matchingBytes_1315(matchingBytes[1315]),
.io_matchingBytes_1316(matchingBytes[1316]),
.io_matchingBytes_1317(matchingBytes[1317]),
.io_matchingBytes_1318(matchingBytes[1318]),
.io_matchingBytes_1319(matchingBytes[1319]),
.io_matchingBytes_1320(matchingBytes[1320]),
.io_matchingBytes_1321(matchingBytes[1321]),
.io_matchingBytes_1322(matchingBytes[1322]),
.io_matchingBytes_1323(matchingBytes[1323]),
.io_matchingBytes_1324(matchingBytes[1324]),
.io_matchingBytes_1325(matchingBytes[1325]),
.io_matchingBytes_1326(matchingBytes[1326]),
.io_matchingBytes_1327(matchingBytes[1327]),
.io_matchingBytes_1328(matchingBytes[1328]),
.io_matchingBytes_1329(matchingBytes[1329]),
.io_matchingBytes_1330(matchingBytes[1330]),
.io_matchingBytes_1331(matchingBytes[1331]),
.io_matchingBytes_1332(matchingBytes[1332]),
.io_matchingBytes_1333(matchingBytes[1333]),
.io_matchingBytes_1334(matchingBytes[1334]),
.io_matchingBytes_1335(matchingBytes[1335]),
.io_matchingBytes_1336(matchingBytes[1336]),
.io_matchingBytes_1337(matchingBytes[1337]),
.io_matchingBytes_1338(matchingBytes[1338]),
.io_matchingBytes_1339(matchingBytes[1339]),
.io_matchingBytes_1340(matchingBytes[1340]),
.io_matchingBytes_1341(matchingBytes[1341]),
.io_matchingBytes_1342(matchingBytes[1342]),
.io_matchingBytes_1343(matchingBytes[1343]),
.io_matchingBytes_1344(matchingBytes[1344]),
.io_matchingBytes_1345(matchingBytes[1345]),
.io_matchingBytes_1346(matchingBytes[1346]),
.io_matchingBytes_1347(matchingBytes[1347]),
.io_matchingBytes_1348(matchingBytes[1348]),
.io_matchingBytes_1349(matchingBytes[1349]),
.io_matchingBytes_1350(matchingBytes[1350]),
.io_matchingBytes_1351(matchingBytes[1351]),
.io_matchingBytes_1352(matchingBytes[1352]),
.io_matchingBytes_1353(matchingBytes[1353]),
.io_matchingBytes_1354(matchingBytes[1354]),
.io_matchingBytes_1355(matchingBytes[1355]),
.io_matchingBytes_1356(matchingBytes[1356]),
.io_matchingBytes_1357(matchingBytes[1357]),
.io_matchingBytes_1358(matchingBytes[1358]),
.io_matchingBytes_1359(matchingBytes[1359]),
.io_matchingBytes_1360(matchingBytes[1360]),
.io_matchingBytes_1361(matchingBytes[1361]),
.io_matchingBytes_1362(matchingBytes[1362]),
.io_matchingBytes_1363(matchingBytes[1363]),
.io_matchingBytes_1364(matchingBytes[1364]),
.io_matchingBytes_1365(matchingBytes[1365]),
.io_matchingBytes_1366(matchingBytes[1366]),
.io_matchingBytes_1367(matchingBytes[1367]),
.io_matchingBytes_1368(matchingBytes[1368]),
.io_matchingBytes_1369(matchingBytes[1369]),
.io_matchingBytes_1370(matchingBytes[1370]),
.io_matchingBytes_1371(matchingBytes[1371]),
.io_matchingBytes_1372(matchingBytes[1372]),
.io_matchingBytes_1373(matchingBytes[1373]),
.io_matchingBytes_1374(matchingBytes[1374]),
.io_matchingBytes_1375(matchingBytes[1375]),
.io_matchingBytes_1376(matchingBytes[1376]),
.io_matchingBytes_1377(matchingBytes[1377]),
.io_matchingBytes_1378(matchingBytes[1378]),
.io_matchingBytes_1379(matchingBytes[1379]),
.io_matchingBytes_1380(matchingBytes[1380]),
.io_matchingBytes_1381(matchingBytes[1381]),
.io_matchingBytes_1382(matchingBytes[1382]),
.io_matchingBytes_1383(matchingBytes[1383]),
.io_matchingBytes_1384(matchingBytes[1384]),
.io_matchingBytes_1385(matchingBytes[1385]),
.io_matchingBytes_1386(matchingBytes[1386]),
.io_matchingBytes_1387(matchingBytes[1387]),
.io_matchingBytes_1388(matchingBytes[1388]),
.io_matchingBytes_1389(matchingBytes[1389]),
.io_matchingBytes_1390(matchingBytes[1390]),
.io_matchingBytes_1391(matchingBytes[1391]),
.io_matchingBytes_1392(matchingBytes[1392]),
.io_matchingBytes_1393(matchingBytes[1393]),
.io_matchingBytes_1394(matchingBytes[1394]),
.io_matchingBytes_1395(matchingBytes[1395]),
.io_matchingBytes_1396(matchingBytes[1396]),
.io_matchingBytes_1397(matchingBytes[1397]),
.io_matchingBytes_1398(matchingBytes[1398]),
.io_matchingBytes_1399(matchingBytes[1399]),
.io_matchingBytes_1400(matchingBytes[1400]),
.io_matchingBytes_1401(matchingBytes[1401]),
.io_matchingBytes_1402(matchingBytes[1402]),
.io_matchingBytes_1403(matchingBytes[1403]),
.io_matchingBytes_1404(matchingBytes[1404]),
.io_matchingBytes_1405(matchingBytes[1405]),
.io_matchingBytes_1406(matchingBytes[1406]),
.io_matchingBytes_1407(matchingBytes[1407]),
.io_matchingBytes_1408(matchingBytes[1408]),
.io_matchingBytes_1409(matchingBytes[1409]),
.io_matchingBytes_1410(matchingBytes[1410]),
.io_matchingBytes_1411(matchingBytes[1411]),
.io_matchingBytes_1412(matchingBytes[1412]),
.io_matchingBytes_1413(matchingBytes[1413]),
.io_matchingBytes_1414(matchingBytes[1414]),
.io_matchingBytes_1415(matchingBytes[1415]),
.io_matchingBytes_1416(matchingBytes[1416]),
.io_matchingBytes_1417(matchingBytes[1417]),
.io_matchingBytes_1418(matchingBytes[1418]),
.io_matchingBytes_1419(matchingBytes[1419]),
.io_matchingBytes_1420(matchingBytes[1420]),
.io_matchingBytes_1421(matchingBytes[1421]),
.io_matchingBytes_1422(matchingBytes[1422]),
.io_matchingBytes_1423(matchingBytes[1423]),
.io_matchingBytes_1424(matchingBytes[1424]),
.io_matchingBytes_1425(matchingBytes[1425]),
.io_matchingBytes_1426(matchingBytes[1426]),
.io_matchingBytes_1427(matchingBytes[1427]),
.io_matchingBytes_1428(matchingBytes[1428]),
.io_matchingBytes_1429(matchingBytes[1429]),
.io_matchingBytes_1430(matchingBytes[1430]),
.io_matchingBytes_1431(matchingBytes[1431]),
.io_matchingBytes_1432(matchingBytes[1432]),
.io_matchingBytes_1433(matchingBytes[1433]),
.io_matchingBytes_1434(matchingBytes[1434]),
.io_matchingBytes_1435(matchingBytes[1435]),
.io_matchingBytes_1436(matchingBytes[1436]),
.io_matchingBytes_1437(matchingBytes[1437]),
.io_matchingBytes_1438(matchingBytes[1438]),
.io_matchingBytes_1439(matchingBytes[1439]),
.io_matchingBytes_1440(matchingBytes[1440]),
.io_matchingBytes_1441(matchingBytes[1441]),
.io_matchingBytes_1442(matchingBytes[1442]),
.io_matchingBytes_1443(matchingBytes[1443]),
.io_matchingBytes_1444(matchingBytes[1444]),
.io_matchingBytes_1445(matchingBytes[1445]),
.io_matchingBytes_1446(matchingBytes[1446]),
.io_matchingBytes_1447(matchingBytes[1447]),
.io_matchingBytes_1448(matchingBytes[1448]),
.io_matchingBytes_1449(matchingBytes[1449]),
.io_matchingBytes_1450(matchingBytes[1450]),
.io_matchingBytes_1451(matchingBytes[1451]),
.io_matchingBytes_1452(matchingBytes[1452]),
.io_matchingBytes_1453(matchingBytes[1453]),
.io_matchingBytes_1454(matchingBytes[1454]),
.io_matchingBytes_1455(matchingBytes[1455]),
.io_matchingBytes_1456(matchingBytes[1456]),
.io_matchingBytes_1457(matchingBytes[1457]),
.io_matchingBytes_1458(matchingBytes[1458]),
.io_matchingBytes_1459(matchingBytes[1459]),
.io_matchingBytes_1460(matchingBytes[1460]),
.io_matchingBytes_1461(matchingBytes[1461]),
.io_matchingBytes_1462(matchingBytes[1462]),
.io_matchingBytes_1463(matchingBytes[1463]),
.io_matchingBytes_1464(matchingBytes[1464]),
.io_matchingBytes_1465(matchingBytes[1465]),
.io_matchingBytes_1466(matchingBytes[1466]),
.io_matchingBytes_1467(matchingBytes[1467]),
.io_matchingBytes_1468(matchingBytes[1468]),
.io_matchingBytes_1469(matchingBytes[1469]),
.io_matchingBytes_1470(matchingBytes[1470]),
.io_matchingBytes_1471(matchingBytes[1471]),
.io_matchingBytes_1472(matchingBytes[1472]),
.io_matchingBytes_1473(matchingBytes[1473]),
.io_matchingBytes_1474(matchingBytes[1474]),
.io_matchingBytes_1475(matchingBytes[1475]),
.io_matchingBytes_1476(matchingBytes[1476]),
.io_matchingBytes_1477(matchingBytes[1477]),
.io_matchingBytes_1478(matchingBytes[1478]),
.io_matchingBytes_1479(matchingBytes[1479]),
.io_matchingBytes_1480(matchingBytes[1480]),
.io_matchingBytes_1481(matchingBytes[1481]),
.io_matchingBytes_1482(matchingBytes[1482]),
.io_matchingBytes_1483(matchingBytes[1483]),
.io_matchingBytes_1484(matchingBytes[1484]),
.io_matchingBytes_1485(matchingBytes[1485]),
.io_matchingBytes_1486(matchingBytes[1486]),
.io_matchingBytes_1487(matchingBytes[1487]),
.io_matchingBytes_1488(matchingBytes[1488]),
.io_matchingBytes_1489(matchingBytes[1489]),
.io_matchingBytes_1490(matchingBytes[1490]),
.io_matchingBytes_1491(matchingBytes[1491]),
.io_matchingBytes_1492(matchingBytes[1492]),
.io_matchingBytes_1493(matchingBytes[1493]),
.io_matchingBytes_1494(matchingBytes[1494]),
.io_matchingBytes_1495(matchingBytes[1495]),
.io_matchingBytes_1496(matchingBytes[1496]),
.io_matchingBytes_1497(matchingBytes[1497]),
.io_matchingBytes_1498(matchingBytes[1498]),
.io_matchingBytes_1499(matchingBytes[1499]),
.io_matchingBytes_1500(matchingBytes[1500]),
.io_matchingBytes_1501(matchingBytes[1501]),
.io_matchingBytes_1502(matchingBytes[1502]),
.io_matchingBytes_1503(matchingBytes[1503]),
.io_matchingBytes_1504(matchingBytes[1504]),
.io_matchingBytes_1505(matchingBytes[1505]),
.io_matchingBytes_1506(matchingBytes[1506]),
.io_matchingBytes_1507(matchingBytes[1507]),
.io_matchingBytes_1508(matchingBytes[1508]),
.io_matchingBytes_1509(matchingBytes[1509]),
.io_matchingBytes_1510(matchingBytes[1510]),
.io_matchingBytes_1511(matchingBytes[1511]),
.io_matchingBytes_1512(matchingBytes[1512]),
.io_matchingBytes_1513(matchingBytes[1513]),
.io_matchingBytes_1514(matchingBytes[1514]),
.io_matchingBytes_1515(matchingBytes[1515]),
.io_matchingBytes_1516(matchingBytes[1516]),
.io_matchingBytes_1517(matchingBytes[1517]),
.io_matchingBytes_1518(matchingBytes[1518]),
.io_matchingBytes_1519(matchingBytes[1519]),
.io_matchingBytes_1520(matchingBytes[1520]),
.io_matchingBytes_1521(matchingBytes[1521]),
.io_matchingBytes_1522(matchingBytes[1522]),
.io_matchingBytes_1523(matchingBytes[1523]),
.io_matchingBytes_1524(matchingBytes[1524]),
.io_matchingBytes_1525(matchingBytes[1525]),
.io_matchingBytes_1526(matchingBytes[1526]),
.io_matchingBytes_1527(matchingBytes[1527]),
.io_matchingBytes_1528(matchingBytes[1528]),
.io_matchingBytes_1529(matchingBytes[1529]),
.io_matchingBytes_1530(matchingBytes[1530]),
.io_matchingBytes_1531(matchingBytes[1531]),
.io_matchingBytes_1532(matchingBytes[1532]),
.io_matchingBytes_1533(matchingBytes[1533]),
.io_matchingBytes_1534(matchingBytes[1534]),
.io_matchingBytes_1535(matchingBytes[1535]),
.io_matchingBytes_1536(matchingBytes[1536]),
.io_matchingBytes_1537(matchingBytes[1537]),
.io_matchingBytes_1538(matchingBytes[1538]),
.io_matchingBytes_1539(matchingBytes[1539]),
.io_matchingBytes_1540(matchingBytes[1540]),
.io_matchingBytes_1541(matchingBytes[1541]),
.io_matchingBytes_1542(matchingBytes[1542]),
.io_matchingBytes_1543(matchingBytes[1543]),
.io_matchingBytes_1544(matchingBytes[1544]),
.io_matchingBytes_1545(matchingBytes[1545]),
.io_matchingBytes_1546(matchingBytes[1546]),
.io_matchingBytes_1547(matchingBytes[1547]),
.io_matchingBytes_1548(matchingBytes[1548]),
.io_matchingBytes_1549(matchingBytes[1549]),
.io_matchingBytes_1550(matchingBytes[1550]),
.io_matchingBytes_1551(matchingBytes[1551]),
.io_matchingBytes_1552(matchingBytes[1552]),
.io_matchingBytes_1553(matchingBytes[1553]),
.io_matchingBytes_1554(matchingBytes[1554]),
.io_matchingBytes_1555(matchingBytes[1555]),
.io_matchingBytes_1556(matchingBytes[1556]),
.io_matchingBytes_1557(matchingBytes[1557]),
.io_matchingBytes_1558(matchingBytes[1558]),
.io_matchingBytes_1559(matchingBytes[1559]),
.io_matchingBytes_1560(matchingBytes[1560]),
.io_matchingBytes_1561(matchingBytes[1561]),
.io_matchingBytes_1562(matchingBytes[1562]),
.io_matchingBytes_1563(matchingBytes[1563]),
.io_matchingBytes_1564(matchingBytes[1564]),
.io_matchingBytes_1565(matchingBytes[1565]),
.io_matchingBytes_1566(matchingBytes[1566]),
.io_matchingBytes_1567(matchingBytes[1567]),
.io_matchingBytes_1568(matchingBytes[1568]),
.io_matchingBytes_1569(matchingBytes[1569]),
.io_matchingBytes_1570(matchingBytes[1570]),
.io_matchingBytes_1571(matchingBytes[1571]),
.io_matchingBytes_1572(matchingBytes[1572]),
.io_matchingBytes_1573(matchingBytes[1573]),
.io_matchingBytes_1574(matchingBytes[1574]),
.io_matchingBytes_1575(matchingBytes[1575]),
.io_matchingBytes_1576(matchingBytes[1576]),
.io_matchingBytes_1577(matchingBytes[1577]),
.io_matchingBytes_1578(matchingBytes[1578]),
.io_matchingBytes_1579(matchingBytes[1579]),
.io_matchingBytes_1580(matchingBytes[1580]),
.io_matchingBytes_1581(matchingBytes[1581]),
.io_matchingBytes_1582(matchingBytes[1582]),
.io_matchingBytes_1583(matchingBytes[1583]),
.io_matchingBytes_1584(matchingBytes[1584]),
.io_matchingBytes_1585(matchingBytes[1585]),
.io_matchingBytes_1586(matchingBytes[1586]),
.io_matchingBytes_1587(matchingBytes[1587]),
.io_matchingBytes_1588(matchingBytes[1588]),
.io_matchingBytes_1589(matchingBytes[1589]),
.io_matchingBytes_1590(matchingBytes[1590]),
.io_matchingBytes_1591(matchingBytes[1591]),
.io_matchingBytes_1592(matchingBytes[1592]),
.io_matchingBytes_1593(matchingBytes[1593]),
.io_matchingBytes_1594(matchingBytes[1594]),
.io_matchingBytes_1595(matchingBytes[1595]),
.io_matchingBytes_1596(matchingBytes[1596]),
.io_matchingBytes_1597(matchingBytes[1597]),
.io_matchingBytes_1598(matchingBytes[1598]),
.io_matchingBytes_1599(matchingBytes[1599]),
.io_matchingBytes_1600(matchingBytes[1600]),
.io_matchingBytes_1601(matchingBytes[1601]),
.io_matchingBytes_1602(matchingBytes[1602]),
.io_matchingBytes_1603(matchingBytes[1603]),
.io_matchingBytes_1604(matchingBytes[1604]),
.io_matchingBytes_1605(matchingBytes[1605]),
.io_matchingBytes_1606(matchingBytes[1606]),
.io_matchingBytes_1607(matchingBytes[1607]),
.io_matchingBytes_1608(matchingBytes[1608]),
.io_matchingBytes_1609(matchingBytes[1609]),
.io_matchingBytes_1610(matchingBytes[1610]),
.io_matchingBytes_1611(matchingBytes[1611]),
.io_matchingBytes_1612(matchingBytes[1612]),
.io_matchingBytes_1613(matchingBytes[1613]),
.io_matchingBytes_1614(matchingBytes[1614]),
.io_matchingBytes_1615(matchingBytes[1615]),
.io_matchingBytes_1616(matchingBytes[1616]),
.io_matchingBytes_1617(matchingBytes[1617]),
.io_matchingBytes_1618(matchingBytes[1618]),
.io_matchingBytes_1619(matchingBytes[1619]),
.io_matchingBytes_1620(matchingBytes[1620]),
.io_matchingBytes_1621(matchingBytes[1621]),
.io_matchingBytes_1622(matchingBytes[1622]),
.io_matchingBytes_1623(matchingBytes[1623]),
.io_matchingBytes_1624(matchingBytes[1624]),
.io_matchingBytes_1625(matchingBytes[1625]),
.io_matchingBytes_1626(matchingBytes[1626]),
.io_matchingBytes_1627(matchingBytes[1627]),
.io_matchingBytes_1628(matchingBytes[1628]),
.io_matchingBytes_1629(matchingBytes[1629]),
.io_matchingBytes_1630(matchingBytes[1630]),
.io_matchingBytes_1631(matchingBytes[1631]),
.io_matchingBytes_1632(matchingBytes[1632]),
.io_matchingBytes_1633(matchingBytes[1633]),
.io_matchingBytes_1634(matchingBytes[1634]),
.io_matchingBytes_1635(matchingBytes[1635]),
.io_matchingBytes_1636(matchingBytes[1636]),
.io_matchingBytes_1637(matchingBytes[1637]),
.io_matchingBytes_1638(matchingBytes[1638]),
.io_matchingBytes_1639(matchingBytes[1639]),
.io_matchingBytes_1640(matchingBytes[1640]),
.io_matchingBytes_1641(matchingBytes[1641]),
.io_matchingBytes_1642(matchingBytes[1642]),
.io_matchingBytes_1643(matchingBytes[1643]),
.io_matchingBytes_1644(matchingBytes[1644]),
.io_matchingBytes_1645(matchingBytes[1645]),
.io_matchingBytes_1646(matchingBytes[1646]),
.io_matchingBytes_1647(matchingBytes[1647]),
.io_matchingBytes_1648(matchingBytes[1648]),
.io_matchingBytes_1649(matchingBytes[1649]),
.io_matchingBytes_1650(matchingBytes[1650]),
.io_matchingBytes_1651(matchingBytes[1651]),
.io_matchingBytes_1652(matchingBytes[1652]),
.io_matchingBytes_1653(matchingBytes[1653]),
.io_matchingBytes_1654(matchingBytes[1654]),
.io_matchingBytes_1655(matchingBytes[1655]),
.io_matchingBytes_1656(matchingBytes[1656]),
.io_matchingBytes_1657(matchingBytes[1657]),
.io_matchingBytes_1658(matchingBytes[1658]),
.io_matchingBytes_1659(matchingBytes[1659]),
.io_matchingBytes_1660(matchingBytes[1660]),
.io_matchingBytes_1661(matchingBytes[1661]),
.io_matchingBytes_1662(matchingBytes[1662]),
.io_matchingBytes_1663(matchingBytes[1663]),
.io_matchingBytes_1664(matchingBytes[1664]),
.io_matchingBytes_1665(matchingBytes[1665]),
.io_matchingBytes_1666(matchingBytes[1666]),
.io_matchingBytes_1667(matchingBytes[1667]),
.io_matchingBytes_1668(matchingBytes[1668]),
.io_matchingBytes_1669(matchingBytes[1669]),
.io_matchingBytes_1670(matchingBytes[1670]),
.io_matchingBytes_1671(matchingBytes[1671]),
.io_matchingBytes_1672(matchingBytes[1672]),
.io_matchingBytes_1673(matchingBytes[1673]),
.io_matchingBytes_1674(matchingBytes[1674]),
.io_matchingBytes_1675(matchingBytes[1675]),
.io_matchingBytes_1676(matchingBytes[1676]),
.io_matchingBytes_1677(matchingBytes[1677]),
.io_matchingBytes_1678(matchingBytes[1678]),
.io_matchingBytes_1679(matchingBytes[1679]),
.io_matchingBytes_1680(matchingBytes[1680]),
.io_matchingBytes_1681(matchingBytes[1681]),
.io_matchingBytes_1682(matchingBytes[1682]),
.io_matchingBytes_1683(matchingBytes[1683]),
.io_matchingBytes_1684(matchingBytes[1684]),
.io_matchingBytes_1685(matchingBytes[1685]),
.io_matchingBytes_1686(matchingBytes[1686]),
.io_matchingBytes_1687(matchingBytes[1687]),
.io_matchingBytes_1688(matchingBytes[1688]),
.io_matchingBytes_1689(matchingBytes[1689]),
.io_matchingBytes_1690(matchingBytes[1690]),
.io_matchingBytes_1691(matchingBytes[1691]),
.io_matchingBytes_1692(matchingBytes[1692]),
.io_matchingBytes_1693(matchingBytes[1693]),
.io_matchingBytes_1694(matchingBytes[1694]),
.io_matchingBytes_1695(matchingBytes[1695]),
.io_matchingBytes_1696(matchingBytes[1696]),
.io_matchingBytes_1697(matchingBytes[1697]),
.io_matchingBytes_1698(matchingBytes[1698]),
.io_matchingBytes_1699(matchingBytes[1699]),
.io_matchingBytes_1700(matchingBytes[1700]),
.io_matchingBytes_1701(matchingBytes[1701]),
.io_matchingBytes_1702(matchingBytes[1702]),
.io_matchingBytes_1703(matchingBytes[1703]),
.io_matchingBytes_1704(matchingBytes[1704]),
.io_matchingBytes_1705(matchingBytes[1705]),
.io_matchingBytes_1706(matchingBytes[1706]),
.io_matchingBytes_1707(matchingBytes[1707]),
.io_matchingBytes_1708(matchingBytes[1708]),
.io_matchingBytes_1709(matchingBytes[1709]),
.io_matchingBytes_1710(matchingBytes[1710]),
.io_matchingBytes_1711(matchingBytes[1711]),
.io_matchingBytes_1712(matchingBytes[1712]),
.io_matchingBytes_1713(matchingBytes[1713]),
.io_matchingBytes_1714(matchingBytes[1714]),
.io_matchingBytes_1715(matchingBytes[1715]),
.io_matchingBytes_1716(matchingBytes[1716]),
.io_matchingBytes_1717(matchingBytes[1717]),
.io_matchingBytes_1718(matchingBytes[1718]),
.io_matchingBytes_1719(matchingBytes[1719]),
.io_matchingBytes_1720(matchingBytes[1720]),
.io_matchingBytes_1721(matchingBytes[1721]),
.io_matchingBytes_1722(matchingBytes[1722]),
.io_matchingBytes_1723(matchingBytes[1723]),
.io_matchingBytes_1724(matchingBytes[1724]),
.io_matchingBytes_1725(matchingBytes[1725]),
.io_matchingBytes_1726(matchingBytes[1726]),
.io_matchingBytes_1727(matchingBytes[1727]),
.io_matchingBytes_1728(matchingBytes[1728]),
.io_matchingBytes_1729(matchingBytes[1729]),
.io_matchingBytes_1730(matchingBytes[1730]),
.io_matchingBytes_1731(matchingBytes[1731]),
.io_matchingBytes_1732(matchingBytes[1732]),
.io_matchingBytes_1733(matchingBytes[1733]),
.io_matchingBytes_1734(matchingBytes[1734]),
.io_matchingBytes_1735(matchingBytes[1735]),
.io_matchingBytes_1736(matchingBytes[1736]),
.io_matchingBytes_1737(matchingBytes[1737]),
.io_matchingBytes_1738(matchingBytes[1738]),
.io_matchingBytes_1739(matchingBytes[1739]),
.io_matchingBytes_1740(matchingBytes[1740]),
.io_matchingBytes_1741(matchingBytes[1741]),
.io_matchingBytes_1742(matchingBytes[1742]),
.io_matchingBytes_1743(matchingBytes[1743]),
.io_matchingBytes_1744(matchingBytes[1744]),
.io_matchingBytes_1745(matchingBytes[1745]),
.io_matchingBytes_1746(matchingBytes[1746]),
.io_matchingBytes_1747(matchingBytes[1747]),
.io_matchingBytes_1748(matchingBytes[1748]),
.io_matchingBytes_1749(matchingBytes[1749]),
.io_matchingBytes_1750(matchingBytes[1750]),
.io_matchingBytes_1751(matchingBytes[1751]),
.io_matchingBytes_1752(matchingBytes[1752]),
.io_matchingBytes_1753(matchingBytes[1753]),
.io_matchingBytes_1754(matchingBytes[1754]),
.io_matchingBytes_1755(matchingBytes[1755]),
.io_matchingBytes_1756(matchingBytes[1756]),
.io_matchingBytes_1757(matchingBytes[1757]),
.io_matchingBytes_1758(matchingBytes[1758]),
.io_matchingBytes_1759(matchingBytes[1759]),
.io_matchingBytes_1760(matchingBytes[1760]),
.io_matchingBytes_1761(matchingBytes[1761]),
.io_matchingBytes_1762(matchingBytes[1762]),
.io_matchingBytes_1763(matchingBytes[1763]),
.io_matchingBytes_1764(matchingBytes[1764]),
.io_matchingBytes_1765(matchingBytes[1765]),
.io_matchingBytes_1766(matchingBytes[1766]),
.io_matchingBytes_1767(matchingBytes[1767]),
.io_matchingBytes_1768(matchingBytes[1768]),
.io_matchingBytes_1769(matchingBytes[1769]),
.io_matchingBytes_1770(matchingBytes[1770]),
.io_matchingBytes_1771(matchingBytes[1771]),
.io_matchingBytes_1772(matchingBytes[1772]),
.io_matchingBytes_1773(matchingBytes[1773]),
.io_matchingBytes_1774(matchingBytes[1774]),
.io_matchingBytes_1775(matchingBytes[1775]),
.io_matchingBytes_1776(matchingBytes[1776]),
.io_matchingBytes_1777(matchingBytes[1777]),
.io_matchingBytes_1778(matchingBytes[1778]),
.io_matchingBytes_1779(matchingBytes[1779]),
.io_matchingBytes_1780(matchingBytes[1780]),
.io_matchingBytes_1781(matchingBytes[1781]),
.io_matchingBytes_1782(matchingBytes[1782]),
.io_matchingBytes_1783(matchingBytes[1783]),
.io_matchingBytes_1784(matchingBytes[1784]),
.io_matchingBytes_1785(matchingBytes[1785]),
.io_matchingBytes_1786(matchingBytes[1786]),
.io_matchingBytes_1787(matchingBytes[1787]),
.io_matchingBytes_1788(matchingBytes[1788]),
.io_matchingBytes_1789(matchingBytes[1789]),
.io_matchingBytes_1790(matchingBytes[1790]),
.io_matchingBytes_1791(matchingBytes[1791]),
.io_matchingBytes_1792(matchingBytes[1792]),
.io_matchingBytes_1793(matchingBytes[1793]),
.io_matchingBytes_1794(matchingBytes[1794]),
.io_matchingBytes_1795(matchingBytes[1795]),
.io_matchingBytes_1796(matchingBytes[1796]),
.io_matchingBytes_1797(matchingBytes[1797]),
.io_matchingBytes_1798(matchingBytes[1798]),
.io_matchingBytes_1799(matchingBytes[1799]),
.io_matchingBytes_1800(matchingBytes[1800]),
.io_matchingBytes_1801(matchingBytes[1801]),
.io_matchingBytes_1802(matchingBytes[1802]),
.io_matchingBytes_1803(matchingBytes[1803]),
.io_matchingBytes_1804(matchingBytes[1804]),
.io_matchingBytes_1805(matchingBytes[1805]),
.io_matchingBytes_1806(matchingBytes[1806]),
.io_matchingBytes_1807(matchingBytes[1807]),
.io_matchingBytes_1808(matchingBytes[1808]),
.io_matchingBytes_1809(matchingBytes[1809]),
.io_matchingBytes_1810(matchingBytes[1810]),
.io_matchingBytes_1811(matchingBytes[1811]),
.io_matchingBytes_1812(matchingBytes[1812]),
.io_matchingBytes_1813(matchingBytes[1813]),
.io_matchingBytes_1814(matchingBytes[1814]),
.io_matchingBytes_1815(matchingBytes[1815]),
.io_matchingBytes_1816(matchingBytes[1816]),
.io_matchingBytes_1817(matchingBytes[1817]),
.io_matchingBytes_1818(matchingBytes[1818]),
.io_matchingBytes_1819(matchingBytes[1819]),
.io_matchingBytes_1820(matchingBytes[1820]),
.io_matchingBytes_1821(matchingBytes[1821]),
.io_matchingBytes_1822(matchingBytes[1822]),
.io_matchingBytes_1823(matchingBytes[1823]),
.io_matchingBytes_1824(matchingBytes[1824]),
.io_matchingBytes_1825(matchingBytes[1825]),
.io_matchingBytes_1826(matchingBytes[1826]),
.io_matchingBytes_1827(matchingBytes[1827]),
.io_matchingBytes_1828(matchingBytes[1828]),
.io_matchingBytes_1829(matchingBytes[1829]),
.io_matchingBytes_1830(matchingBytes[1830]),
.io_matchingBytes_1831(matchingBytes[1831]),
.io_matchingBytes_1832(matchingBytes[1832]),
.io_matchingBytes_1833(matchingBytes[1833]),
.io_matchingBytes_1834(matchingBytes[1834]),
.io_matchingBytes_1835(matchingBytes[1835]),
.io_matchingBytes_1836(matchingBytes[1836]),
.io_matchingBytes_1837(matchingBytes[1837]),
.io_matchingBytes_1838(matchingBytes[1838]),
.io_matchingBytes_1839(matchingBytes[1839]),
.io_matchingBytes_1840(matchingBytes[1840]),
.io_matchingBytes_1841(matchingBytes[1841]),
.io_matchingBytes_1842(matchingBytes[1842]),
.io_matchingBytes_1843(matchingBytes[1843]),
.io_matchingBytes_1844(matchingBytes[1844]),
.io_matchingBytes_1845(matchingBytes[1845]),
.io_matchingBytes_1846(matchingBytes[1846]),
.io_matchingBytes_1847(matchingBytes[1847]),
.io_matchingBytes_1848(matchingBytes[1848]),
.io_matchingBytes_1849(matchingBytes[1849]),
.io_matchingBytes_1850(matchingBytes[1850]),
.io_matchingBytes_1851(matchingBytes[1851]),
.io_matchingBytes_1852(matchingBytes[1852]),
.io_matchingBytes_1853(matchingBytes[1853]),
.io_matchingBytes_1854(matchingBytes[1854]),
.io_matchingBytes_1855(matchingBytes[1855]),
.io_matchingBytes_1856(matchingBytes[1856]),
.io_matchingBytes_1857(matchingBytes[1857]),
.io_matchingBytes_1858(matchingBytes[1858]),
.io_matchingBytes_1859(matchingBytes[1859]),
.io_matchingBytes_1860(matchingBytes[1860]),
.io_matchingBytes_1861(matchingBytes[1861]),
.io_matchingBytes_1862(matchingBytes[1862]),
.io_matchingBytes_1863(matchingBytes[1863]),
.io_matchingBytes_1864(matchingBytes[1864]),
.io_matchingBytes_1865(matchingBytes[1865]),
.io_matchingBytes_1866(matchingBytes[1866]),
.io_matchingBytes_1867(matchingBytes[1867]),
.io_matchingBytes_1868(matchingBytes[1868]),
.io_matchingBytes_1869(matchingBytes[1869]),
.io_matchingBytes_1870(matchingBytes[1870]),
.io_matchingBytes_1871(matchingBytes[1871]),
.io_matchingBytes_1872(matchingBytes[1872]),
.io_matchingBytes_1873(matchingBytes[1873]),
.io_matchingBytes_1874(matchingBytes[1874]),
.io_matchingBytes_1875(matchingBytes[1875]),
.io_matchingBytes_1876(matchingBytes[1876]),
.io_matchingBytes_1877(matchingBytes[1877]),
.io_matchingBytes_1878(matchingBytes[1878]),
.io_matchingBytes_1879(matchingBytes[1879]),
.io_matchingBytes_1880(matchingBytes[1880]),
.io_matchingBytes_1881(matchingBytes[1881]),
.io_matchingBytes_1882(matchingBytes[1882]),
.io_matchingBytes_1883(matchingBytes[1883]),
.io_matchingBytes_1884(matchingBytes[1884]),
.io_matchingBytes_1885(matchingBytes[1885]),
.io_matchingBytes_1886(matchingBytes[1886]),
.io_matchingBytes_1887(matchingBytes[1887]),
.io_matchingBytes_1888(matchingBytes[1888]),
.io_matchingBytes_1889(matchingBytes[1889]),
.io_matchingBytes_1890(matchingBytes[1890]),
.io_matchingBytes_1891(matchingBytes[1891]),
.io_matchingBytes_1892(matchingBytes[1892]),
.io_matchingBytes_1893(matchingBytes[1893]),
.io_matchingBytes_1894(matchingBytes[1894]),
.io_matchingBytes_1895(matchingBytes[1895]),
.io_matchingBytes_1896(matchingBytes[1896]),
.io_matchingBytes_1897(matchingBytes[1897]),
.io_matchingBytes_1898(matchingBytes[1898]),
.io_matchingBytes_1899(matchingBytes[1899]),
.io_matchingBytes_1900(matchingBytes[1900]),
.io_matchingBytes_1901(matchingBytes[1901]),
.io_matchingBytes_1902(matchingBytes[1902]),
.io_matchingBytes_1903(matchingBytes[1903]),
.io_matchingBytes_1904(matchingBytes[1904]),
.io_matchingBytes_1905(matchingBytes[1905]),
.io_matchingBytes_1906(matchingBytes[1906]),
.io_matchingBytes_1907(matchingBytes[1907]),
.io_matchingBytes_1908(matchingBytes[1908]),
.io_matchingBytes_1909(matchingBytes[1909]),
.io_matchingBytes_1910(matchingBytes[1910]),
.io_matchingBytes_1911(matchingBytes[1911]),
.io_matchingBytes_1912(matchingBytes[1912]),
.io_matchingBytes_1913(matchingBytes[1913]),
.io_matchingBytes_1914(matchingBytes[1914]),
.io_matchingBytes_1915(matchingBytes[1915]),
.io_matchingBytes_1916(matchingBytes[1916]),
.io_matchingBytes_1917(matchingBytes[1917]),
.io_matchingBytes_1918(matchingBytes[1918]),
.io_matchingBytes_1919(matchingBytes[1919]),
.io_matchingBytes_1920(matchingBytes[1920]),
.io_matchingBytes_1921(matchingBytes[1921]),
.io_matchingBytes_1922(matchingBytes[1922]),
.io_matchingBytes_1923(matchingBytes[1923]),
.io_matchingBytes_1924(matchingBytes[1924]),
.io_matchingBytes_1925(matchingBytes[1925]),
.io_matchingBytes_1926(matchingBytes[1926]),
.io_matchingBytes_1927(matchingBytes[1927]),
.io_matchingBytes_1928(matchingBytes[1928]),
.io_matchingBytes_1929(matchingBytes[1929]),
.io_matchingBytes_1930(matchingBytes[1930]),
.io_matchingBytes_1931(matchingBytes[1931]),
.io_matchingBytes_1932(matchingBytes[1932]),
.io_matchingBytes_1933(matchingBytes[1933]),
.io_matchingBytes_1934(matchingBytes[1934]),
.io_matchingBytes_1935(matchingBytes[1935]),
.io_matchingBytes_1936(matchingBytes[1936]),
.io_matchingBytes_1937(matchingBytes[1937]),
.io_matchingBytes_1938(matchingBytes[1938]),
.io_matchingBytes_1939(matchingBytes[1939]),
.io_matchingBytes_1940(matchingBytes[1940]),
.io_matchingBytes_1941(matchingBytes[1941]),
.io_matchingBytes_1942(matchingBytes[1942]),
.io_matchingBytes_1943(matchingBytes[1943]),
.io_matchingBytes_1944(matchingBytes[1944]),
.io_matchingBytes_1945(matchingBytes[1945]),
.io_matchingBytes_1946(matchingBytes[1946]),
.io_matchingBytes_1947(matchingBytes[1947]),
.io_matchingBytes_1948(matchingBytes[1948]),
.io_matchingBytes_1949(matchingBytes[1949]),
.io_matchingBytes_1950(matchingBytes[1950]),
.io_matchingBytes_1951(matchingBytes[1951]),
.io_matchingBytes_1952(matchingBytes[1952]),
.io_matchingBytes_1953(matchingBytes[1953]),
.io_matchingBytes_1954(matchingBytes[1954]),
.io_matchingBytes_1955(matchingBytes[1955]),
.io_matchingBytes_1956(matchingBytes[1956]),
.io_matchingBytes_1957(matchingBytes[1957]),
.io_matchingBytes_1958(matchingBytes[1958]),
.io_matchingBytes_1959(matchingBytes[1959]),
.io_matchingBytes_1960(matchingBytes[1960]),
.io_matchingBytes_1961(matchingBytes[1961]),
.io_matchingBytes_1962(matchingBytes[1962]),
.io_matchingBytes_1963(matchingBytes[1963]),
.io_matchingBytes_1964(matchingBytes[1964]),
.io_matchingBytes_1965(matchingBytes[1965]),
.io_matchingBytes_1966(matchingBytes[1966]),
.io_matchingBytes_1967(matchingBytes[1967]),
.io_matchingBytes_1968(matchingBytes[1968]),
.io_matchingBytes_1969(matchingBytes[1969]),
.io_matchingBytes_1970(matchingBytes[1970]),
.io_matchingBytes_1971(matchingBytes[1971]),
.io_matchingBytes_1972(matchingBytes[1972]),
.io_matchingBytes_1973(matchingBytes[1973]),
.io_matchingBytes_1974(matchingBytes[1974]),
.io_matchingBytes_1975(matchingBytes[1975]),
.io_matchingBytes_1976(matchingBytes[1976]),
.io_matchingBytes_1977(matchingBytes[1977]),
.io_matchingBytes_1978(matchingBytes[1978]),
.io_matchingBytes_1979(matchingBytes[1979]),
.io_matchingBytes_1980(matchingBytes[1980]),
.io_matchingBytes_1981(matchingBytes[1981]),
.io_matchingBytes_1982(matchingBytes[1982]),
.io_matchingBytes_1983(matchingBytes[1983]),
.io_matchingBytes_1984(matchingBytes[1984]),
.io_matchingBytes_1985(matchingBytes[1985]),
.io_matchingBytes_1986(matchingBytes[1986]),
.io_matchingBytes_1987(matchingBytes[1987]),
.io_matchingBytes_1988(matchingBytes[1988]),
.io_matchingBytes_1989(matchingBytes[1989]),
.io_matchingBytes_1990(matchingBytes[1990]),
.io_matchingBytes_1991(matchingBytes[1991]),
.io_matchingBytes_1992(matchingBytes[1992]),
.io_matchingBytes_1993(matchingBytes[1993]),
.io_matchingBytes_1994(matchingBytes[1994]),
.io_matchingBytes_1995(matchingBytes[1995]),
.io_matchingBytes_1996(matchingBytes[1996]),
.io_matchingBytes_1997(matchingBytes[1997]),
.io_matchingBytes_1998(matchingBytes[1998]),
.io_matchingBytes_1999(matchingBytes[1999]),
.io_matchingBytes_2000(matchingBytes[2000]),
.io_matchingBytes_2001(matchingBytes[2001]),
.io_matchingBytes_2002(matchingBytes[2002]),
.io_matchingBytes_2003(matchingBytes[2003]),
.io_matchingBytes_2004(matchingBytes[2004]),
.io_matchingBytes_2005(matchingBytes[2005]),
.io_matchingBytes_2006(matchingBytes[2006]),
.io_matchingBytes_2007(matchingBytes[2007]),
.io_matchingBytes_2008(matchingBytes[2008]),
.io_matchingBytes_2009(matchingBytes[2009]),
.io_matchingBytes_2010(matchingBytes[2010]),
.io_matchingBytes_2011(matchingBytes[2011]),
.io_matchingBytes_2012(matchingBytes[2012]),
.io_matchingBytes_2013(matchingBytes[2013]),
.io_matchingBytes_2014(matchingBytes[2014]),
.io_matchingBytes_2015(matchingBytes[2015]),
.io_matchingBytes_2016(matchingBytes[2016]),
.io_matchingBytes_2017(matchingBytes[2017]),
.io_matchingBytes_2018(matchingBytes[2018]),
.io_matchingBytes_2019(matchingBytes[2019]),
.io_matchingBytes_2020(matchingBytes[2020]),
.io_matchingBytes_2021(matchingBytes[2021]),
.io_matchingBytes_2022(matchingBytes[2022]),
.io_matchingBytes_2023(matchingBytes[2023]),
.io_matchingBytes_2024(matchingBytes[2024]),
.io_matchingBytes_2025(matchingBytes[2025]),
.io_matchingBytes_2026(matchingBytes[2026]),
.io_matchingBytes_2027(matchingBytes[2027]),
.io_matchingBytes_2028(matchingBytes[2028]),
.io_matchingBytes_2029(matchingBytes[2029]),
.io_matchingBytes_2030(matchingBytes[2030]),
.io_matchingBytes_2031(matchingBytes[2031]),
.io_matchingBytes_2032(matchingBytes[2032]),
.io_matchingBytes_2033(matchingBytes[2033]),
.io_matchingBytes_2034(matchingBytes[2034]),
.io_matchingBytes_2035(matchingBytes[2035]),
.io_matchingBytes_2036(matchingBytes[2036]),
.io_matchingBytes_2037(matchingBytes[2037]),
.io_matchingBytes_2038(matchingBytes[2038]),
.io_matchingBytes_2039(matchingBytes[2039]),
.io_matchingBytes_2040(matchingBytes[2040]),
.io_matchingBytes_2041(matchingBytes[2041]),
.io_matchingBytes_2042(matchingBytes[2042]),
.io_matchingBytes_2043(matchingBytes[2043]),
.io_matchingBytes_2044(matchingBytes[2044]),
.io_matchingBytes_2045(matchingBytes[2045]),
.io_matchingBytes_2046(matchingBytes[2046]),
.io_matchingBytes_2047(matchingBytes[2047]),
.io_matchingBytes_2048(matchingBytes[2048]),
.io_matchingBytes_2049(matchingBytes[2049]),
.io_matchingBytes_2050(matchingBytes[2050]),
.io_matchingBytes_2051(matchingBytes[2051]),
.io_matchingBytes_2052(matchingBytes[2052]),
.io_matchingBytes_2053(matchingBytes[2053]),
.io_matchingBytes_2054(matchingBytes[2054]),
.io_matchingBytes_2055(matchingBytes[2055]),
.io_matchingBytes_2056(matchingBytes[2056]),
.io_matchingBytes_2057(matchingBytes[2057]),
.io_matchingBytes_2058(matchingBytes[2058]),
.io_matchingBytes_2059(matchingBytes[2059]),
.io_matchingBytes_2060(matchingBytes[2060]),
.io_matchingBytes_2061(matchingBytes[2061]),
.io_matchingBytes_2062(matchingBytes[2062]),
.io_matchingBytes_2063(matchingBytes[2063]),
.io_matchingBytes_2064(matchingBytes[2064]),
.io_matchingBytes_2065(matchingBytes[2065]),
.io_matchingBytes_2066(matchingBytes[2066]),
.io_matchingBytes_2067(matchingBytes[2067]),
.io_matchingBytes_2068(matchingBytes[2068]),
.io_matchingBytes_2069(matchingBytes[2069]),
.io_matchingBytes_2070(matchingBytes[2070]),
.io_matchingBytes_2071(matchingBytes[2071]),
.io_matchingBytes_2072(matchingBytes[2072]),
.io_matchingBytes_2073(matchingBytes[2073]),
.io_matchingBytes_2074(matchingBytes[2074]),
.io_matchingBytes_2075(matchingBytes[2075]),
.io_matchingBytes_2076(matchingBytes[2076]),
.io_matchingBytes_2077(matchingBytes[2077]),
.io_matchingBytes_2078(matchingBytes[2078]),
.io_matchingBytes_2079(matchingBytes[2079]),
.io_matchingBytes_2080(matchingBytes[2080]),
.io_matchingBytes_2081(matchingBytes[2081]),
.io_matchingBytes_2082(matchingBytes[2082]),
.io_matchingBytes_2083(matchingBytes[2083]),
.io_matchingBytes_2084(matchingBytes[2084]),
.io_matchingBytes_2085(matchingBytes[2085]),
.io_matchingBytes_2086(matchingBytes[2086]),
.io_matchingBytes_2087(matchingBytes[2087]),
.io_matchingBytes_2088(matchingBytes[2088]),
.io_matchingBytes_2089(matchingBytes[2089]),
.io_matchingBytes_2090(matchingBytes[2090]),
.io_matchingBytes_2091(matchingBytes[2091]),
.io_matchingBytes_2092(matchingBytes[2092]),
.io_matchingBytes_2093(matchingBytes[2093]),
.io_matchingBytes_2094(matchingBytes[2094]),
.io_matchingBytes_2095(matchingBytes[2095]),
.io_matchingBytes_2096(matchingBytes[2096]),
.io_matchingBytes_2097(matchingBytes[2097]),
.io_matchingBytes_2098(matchingBytes[2098]),
.io_matchingBytes_2099(matchingBytes[2099]),
.io_matchingBytes_2100(matchingBytes[2100]),
.io_matchingBytes_2101(matchingBytes[2101]),
.io_matchingBytes_2102(matchingBytes[2102]),
.io_matchingBytes_2103(matchingBytes[2103]),
.io_matchingBytes_2104(matchingBytes[2104]),
.io_matchingBytes_2105(matchingBytes[2105]),
.io_matchingBytes_2106(matchingBytes[2106]),
.io_matchingBytes_2107(matchingBytes[2107]),
.io_matchingBytes_2108(matchingBytes[2108]),
.io_matchingBytes_2109(matchingBytes[2109]),
.io_matchingBytes_2110(matchingBytes[2110]),
.io_matchingBytes_2111(matchingBytes[2111]),
.io_matchingBytes_2112(matchingBytes[2112]),
.io_matchingBytes_2113(matchingBytes[2113]),
.io_matchingBytes_2114(matchingBytes[2114]),
.io_matchingBytes_2115(matchingBytes[2115]),
.io_matchingBytes_2116(matchingBytes[2116]),
.io_matchingBytes_2117(matchingBytes[2117]),
.io_matchingBytes_2118(matchingBytes[2118]),
.io_matchingBytes_2119(matchingBytes[2119]),
.io_matchingBytes_2120(matchingBytes[2120]),
.io_matchingBytes_2121(matchingBytes[2121]),
.io_matchingBytes_2122(matchingBytes[2122]),
.io_matchingBytes_2123(matchingBytes[2123]),
.io_matchingBytes_2124(matchingBytes[2124]),
.io_matchingBytes_2125(matchingBytes[2125]),
.io_matchingBytes_2126(matchingBytes[2126]),
.io_matchingBytes_2127(matchingBytes[2127]),
.io_matchingBytes_2128(matchingBytes[2128]),
.io_matchingBytes_2129(matchingBytes[2129]),
.io_matchingBytes_2130(matchingBytes[2130]),
.io_matchingBytes_2131(matchingBytes[2131]),
.io_matchingBytes_2132(matchingBytes[2132]),
.io_matchingBytes_2133(matchingBytes[2133]),
.io_matchingBytes_2134(matchingBytes[2134]),
.io_matchingBytes_2135(matchingBytes[2135]),
.io_matchingBytes_2136(matchingBytes[2136]),
.io_matchingBytes_2137(matchingBytes[2137]),
.io_matchingBytes_2138(matchingBytes[2138]),
.io_matchingBytes_2139(matchingBytes[2139]),
.io_matchingBytes_2140(matchingBytes[2140]),
.io_matchingBytes_2141(matchingBytes[2141]),
.io_matchingBytes_2142(matchingBytes[2142]),
.io_matchingBytes_2143(matchingBytes[2143]),
.io_matchingBytes_2144(matchingBytes[2144]),
.io_matchingBytes_2145(matchingBytes[2145]),
.io_matchingBytes_2146(matchingBytes[2146]),
.io_matchingBytes_2147(matchingBytes[2147]),
.io_matchingBytes_2148(matchingBytes[2148]),
.io_matchingBytes_2149(matchingBytes[2149]),
.io_matchingBytes_2150(matchingBytes[2150]),
.io_matchingBytes_2151(matchingBytes[2151]),
.io_matchingBytes_2152(matchingBytes[2152]),
.io_matchingBytes_2153(matchingBytes[2153]),
.io_matchingBytes_2154(matchingBytes[2154]),
.io_matchingBytes_2155(matchingBytes[2155]),
.io_matchingBytes_2156(matchingBytes[2156]),
.io_matchingBytes_2157(matchingBytes[2157]),
.io_matchingBytes_2158(matchingBytes[2158]),
.io_matchingBytes_2159(matchingBytes[2159]),
.io_matchingBytes_2160(matchingBytes[2160]),
.io_matchingBytes_2161(matchingBytes[2161]),
.io_matchingBytes_2162(matchingBytes[2162]),
.io_matchingBytes_2163(matchingBytes[2163]),
.io_matchingBytes_2164(matchingBytes[2164]),
.io_matchingBytes_2165(matchingBytes[2165]),
.io_matchingBytes_2166(matchingBytes[2166]),
.io_matchingBytes_2167(matchingBytes[2167]),
.io_matchingBytes_2168(matchingBytes[2168]),
.io_matchingBytes_2169(matchingBytes[2169]),
.io_matchingBytes_2170(matchingBytes[2170]),
.io_matchingBytes_2171(matchingBytes[2171]),
.io_matchingBytes_2172(matchingBytes[2172]),
.io_matchingBytes_2173(matchingBytes[2173]),
.io_matchingBytes_2174(matchingBytes[2174]),
.io_matchingBytes_2175(matchingBytes[2175]),
.io_matchingBytes_2176(matchingBytes[2176]),
.io_matchingBytes_2177(matchingBytes[2177]),
.io_matchingBytes_2178(matchingBytes[2178]),
.io_matchingBytes_2179(matchingBytes[2179]),
.io_matchingBytes_2180(matchingBytes[2180]),
.io_matchingBytes_2181(matchingBytes[2181]),
.io_matchingBytes_2182(matchingBytes[2182]),
.io_matchingBytes_2183(matchingBytes[2183]),
.io_matchingBytes_2184(matchingBytes[2184]),
.io_matchingBytes_2185(matchingBytes[2185]),
.io_matchingBytes_2186(matchingBytes[2186]),
.io_matchingBytes_2187(matchingBytes[2187]),
.io_matchingBytes_2188(matchingBytes[2188]),
.io_matchingBytes_2189(matchingBytes[2189]),
.io_matchingBytes_2190(matchingBytes[2190]),
.io_matchingBytes_2191(matchingBytes[2191]),
.io_matchingBytes_2192(matchingBytes[2192]),
.io_matchingBytes_2193(matchingBytes[2193]),
.io_matchingBytes_2194(matchingBytes[2194]),
.io_matchingBytes_2195(matchingBytes[2195]),
.io_matchingBytes_2196(matchingBytes[2196]),
.io_matchingBytes_2197(matchingBytes[2197]),
.io_matchingBytes_2198(matchingBytes[2198]),
.io_matchingBytes_2199(matchingBytes[2199]),
.io_matchingBytes_2200(matchingBytes[2200]),
.io_matchingBytes_2201(matchingBytes[2201]),
.io_matchingBytes_2202(matchingBytes[2202]),
.io_matchingBytes_2203(matchingBytes[2203]),
.io_matchingBytes_2204(matchingBytes[2204]),
.io_matchingBytes_2205(matchingBytes[2205]),
.io_matchingBytes_2206(matchingBytes[2206]),
.io_matchingBytes_2207(matchingBytes[2207]),
.io_matchingBytes_2208(matchingBytes[2208]),
.io_matchingBytes_2209(matchingBytes[2209]),
.io_matchingBytes_2210(matchingBytes[2210]),
.io_matchingBytes_2211(matchingBytes[2211]),
.io_matchingBytes_2212(matchingBytes[2212]),
.io_matchingBytes_2213(matchingBytes[2213]),
.io_matchingBytes_2214(matchingBytes[2214]),
.io_matchingBytes_2215(matchingBytes[2215]),
.io_matchingBytes_2216(matchingBytes[2216]),
.io_matchingBytes_2217(matchingBytes[2217]),
.io_matchingBytes_2218(matchingBytes[2218]),
.io_matchingBytes_2219(matchingBytes[2219]),
.io_matchingBytes_2220(matchingBytes[2220]),
.io_matchingBytes_2221(matchingBytes[2221]),
.io_matchingBytes_2222(matchingBytes[2222]),
.io_matchingBytes_2223(matchingBytes[2223]),
.io_matchingBytes_2224(matchingBytes[2224]),
.io_matchingBytes_2225(matchingBytes[2225]),
.io_matchingBytes_2226(matchingBytes[2226]),
.io_matchingBytes_2227(matchingBytes[2227]),
.io_matchingBytes_2228(matchingBytes[2228]),
.io_matchingBytes_2229(matchingBytes[2229]),
.io_matchingBytes_2230(matchingBytes[2230]),
.io_matchingBytes_2231(matchingBytes[2231]),
.io_matchingBytes_2232(matchingBytes[2232]),
.io_matchingBytes_2233(matchingBytes[2233]),
.io_matchingBytes_2234(matchingBytes[2234]),
.io_matchingBytes_2235(matchingBytes[2235]),
.io_matchingBytes_2236(matchingBytes[2236]),
.io_matchingBytes_2237(matchingBytes[2237]),
.io_matchingBytes_2238(matchingBytes[2238]),
.io_matchingBytes_2239(matchingBytes[2239]),
.io_matchingBytes_2240(matchingBytes[2240]),
.io_matchingBytes_2241(matchingBytes[2241]),
.io_matchingBytes_2242(matchingBytes[2242]),
.io_matchingBytes_2243(matchingBytes[2243]),
.io_matchingBytes_2244(matchingBytes[2244]),
.io_matchingBytes_2245(matchingBytes[2245]),
.io_matchingBytes_2246(matchingBytes[2246]),
.io_matchingBytes_2247(matchingBytes[2247]),
.io_matchingBytes_2248(matchingBytes[2248]),
.io_matchingBytes_2249(matchingBytes[2249]),
.io_matchingBytes_2250(matchingBytes[2250]),
.io_matchingBytes_2251(matchingBytes[2251]),
.io_matchingBytes_2252(matchingBytes[2252]),
.io_matchingBytes_2253(matchingBytes[2253]),
.io_matchingBytes_2254(matchingBytes[2254]),
.io_matchingBytes_2255(matchingBytes[2255]),
.io_matchingBytes_2256(matchingBytes[2256]),
.io_matchingBytes_2257(matchingBytes[2257]),
.io_matchingBytes_2258(matchingBytes[2258]),
.io_matchingBytes_2259(matchingBytes[2259]),
.io_matchingBytes_2260(matchingBytes[2260]),
.io_matchingBytes_2261(matchingBytes[2261]),
.io_matchingBytes_2262(matchingBytes[2262]),
.io_matchingBytes_2263(matchingBytes[2263]),
.io_matchingBytes_2264(matchingBytes[2264]),
.io_matchingBytes_2265(matchingBytes[2265]),
.io_matchingBytes_2266(matchingBytes[2266]),
.io_matchingBytes_2267(matchingBytes[2267]),
.io_matchingBytes_2268(matchingBytes[2268]),
.io_matchingBytes_2269(matchingBytes[2269]),
.io_matchingBytes_2270(matchingBytes[2270]),
.io_matchingBytes_2271(matchingBytes[2271]),
.io_matchingBytes_2272(matchingBytes[2272]),
.io_matchingBytes_2273(matchingBytes[2273]),
.io_matchingBytes_2274(matchingBytes[2274]),
.io_matchingBytes_2275(matchingBytes[2275]),
.io_matchingBytes_2276(matchingBytes[2276]),
.io_matchingBytes_2277(matchingBytes[2277]),
.io_matchingBytes_2278(matchingBytes[2278]),
.io_matchingBytes_2279(matchingBytes[2279]),
.io_matchingBytes_2280(matchingBytes[2280]),
.io_matchingBytes_2281(matchingBytes[2281]),
.io_matchingBytes_2282(matchingBytes[2282]),
.io_matchingBytes_2283(matchingBytes[2283]),
.io_matchingBytes_2284(matchingBytes[2284]),
.io_matchingBytes_2285(matchingBytes[2285]),
.io_matchingBytes_2286(matchingBytes[2286]),
.io_matchingBytes_2287(matchingBytes[2287]),
.io_matchingBytes_2288(matchingBytes[2288]),
.io_matchingBytes_2289(matchingBytes[2289]),
.io_matchingBytes_2290(matchingBytes[2290]),
.io_matchingBytes_2291(matchingBytes[2291]),
.io_matchingBytes_2292(matchingBytes[2292]),
.io_matchingBytes_2293(matchingBytes[2293]),
.io_matchingBytes_2294(matchingBytes[2294]),
.io_matchingBytes_2295(matchingBytes[2295]),
.io_matchingBytes_2296(matchingBytes[2296]),
.io_matchingBytes_2297(matchingBytes[2297]),
.io_matchingBytes_2298(matchingBytes[2298]),
.io_matchingBytes_2299(matchingBytes[2299]),
.io_matchingBytes_2300(matchingBytes[2300]),
.io_matchingBytes_2301(matchingBytes[2301]),
.io_matchingBytes_2302(matchingBytes[2302]),
.io_matchingBytes_2303(matchingBytes[2303]),
.io_matchingBytes_2304(matchingBytes[2304]),
.io_matchingBytes_2305(matchingBytes[2305]),
.io_matchingBytes_2306(matchingBytes[2306]),
.io_matchingBytes_2307(matchingBytes[2307]),
.io_matchingBytes_2308(matchingBytes[2308]),
.io_matchingBytes_2309(matchingBytes[2309]),
.io_matchingBytes_2310(matchingBytes[2310]),
.io_matchingBytes_2311(matchingBytes[2311]),
.io_matchingBytes_2312(matchingBytes[2312]),
.io_matchingBytes_2313(matchingBytes[2313]),
.io_matchingBytes_2314(matchingBytes[2314]),
.io_matchingBytes_2315(matchingBytes[2315]),
.io_matchingBytes_2316(matchingBytes[2316]),
.io_matchingBytes_2317(matchingBytes[2317]),
.io_matchingBytes_2318(matchingBytes[2318]),
.io_matchingBytes_2319(matchingBytes[2319]),
.io_matchingBytes_2320(matchingBytes[2320]),
.io_matchingBytes_2321(matchingBytes[2321]),
.io_matchingBytes_2322(matchingBytes[2322]),
.io_matchingBytes_2323(matchingBytes[2323]),
.io_matchingBytes_2324(matchingBytes[2324]),
.io_matchingBytes_2325(matchingBytes[2325]),
.io_matchingBytes_2326(matchingBytes[2326]),
.io_matchingBytes_2327(matchingBytes[2327]),
.io_matchingBytes_2328(matchingBytes[2328]),
.io_matchingBytes_2329(matchingBytes[2329]),
.io_matchingBytes_2330(matchingBytes[2330]),
.io_matchingBytes_2331(matchingBytes[2331]),
.io_matchingBytes_2332(matchingBytes[2332]),
.io_matchingBytes_2333(matchingBytes[2333]),
.io_matchingBytes_2334(matchingBytes[2334]),
.io_matchingBytes_2335(matchingBytes[2335]),
.io_matchingBytes_2336(matchingBytes[2336]),
.io_matchingBytes_2337(matchingBytes[2337]),
.io_matchingBytes_2338(matchingBytes[2338]),
.io_matchingBytes_2339(matchingBytes[2339]),
.io_matchingBytes_2340(matchingBytes[2340]),
.io_matchingBytes_2341(matchingBytes[2341]),
.io_matchingBytes_2342(matchingBytes[2342]),
.io_matchingBytes_2343(matchingBytes[2343]),
.io_matchingBytes_2344(matchingBytes[2344]),
.io_matchingBytes_2345(matchingBytes[2345]),
.io_matchingBytes_2346(matchingBytes[2346]),
.io_matchingBytes_2347(matchingBytes[2347]),
.io_matchingBytes_2348(matchingBytes[2348]),
.io_matchingBytes_2349(matchingBytes[2349]),
.io_matchingBytes_2350(matchingBytes[2350]),
.io_matchingBytes_2351(matchingBytes[2351]),
.io_matchingBytes_2352(matchingBytes[2352]),
.io_matchingBytes_2353(matchingBytes[2353]),
.io_matchingBytes_2354(matchingBytes[2354]),
.io_matchingBytes_2355(matchingBytes[2355]),
.io_matchingBytes_2356(matchingBytes[2356]),
.io_matchingBytes_2357(matchingBytes[2357]),
.io_matchingBytes_2358(matchingBytes[2358]),
.io_matchingBytes_2359(matchingBytes[2359]),
.io_matchingBytes_2360(matchingBytes[2360]),
.io_matchingBytes_2361(matchingBytes[2361]),
.io_matchingBytes_2362(matchingBytes[2362]),
.io_matchingBytes_2363(matchingBytes[2363]),
.io_matchingBytes_2364(matchingBytes[2364]),
.io_matchingBytes_2365(matchingBytes[2365]),
.io_matchingBytes_2366(matchingBytes[2366]),
.io_matchingBytes_2367(matchingBytes[2367]),
.io_matchingBytes_2368(matchingBytes[2368]),
.io_matchingBytes_2369(matchingBytes[2369]),
.io_matchingBytes_2370(matchingBytes[2370]),
.io_matchingBytes_2371(matchingBytes[2371]),
.io_matchingBytes_2372(matchingBytes[2372]),
.io_matchingBytes_2373(matchingBytes[2373]),
.io_matchingBytes_2374(matchingBytes[2374]),
.io_matchingBytes_2375(matchingBytes[2375]),
.io_matchingBytes_2376(matchingBytes[2376]),
.io_matchingBytes_2377(matchingBytes[2377]),
.io_matchingBytes_2378(matchingBytes[2378]),
.io_matchingBytes_2379(matchingBytes[2379]),
.io_matchingBytes_2380(matchingBytes[2380]),
.io_matchingBytes_2381(matchingBytes[2381]),
.io_matchingBytes_2382(matchingBytes[2382]),
.io_matchingBytes_2383(matchingBytes[2383]),
.io_matchingBytes_2384(matchingBytes[2384]),
.io_matchingBytes_2385(matchingBytes[2385]),
.io_matchingBytes_2386(matchingBytes[2386]),
.io_matchingBytes_2387(matchingBytes[2387]),
.io_matchingBytes_2388(matchingBytes[2388]),
.io_matchingBytes_2389(matchingBytes[2389]),
.io_matchingBytes_2390(matchingBytes[2390]),
.io_matchingBytes_2391(matchingBytes[2391]),
.io_matchingBytes_2392(matchingBytes[2392]),
.io_matchingBytes_2393(matchingBytes[2393]),
.io_matchingBytes_2394(matchingBytes[2394]),
.io_matchingBytes_2395(matchingBytes[2395]),
.io_matchingBytes_2396(matchingBytes[2396]),
.io_matchingBytes_2397(matchingBytes[2397]),
.io_matchingBytes_2398(matchingBytes[2398]),
.io_matchingBytes_2399(matchingBytes[2399]),
.io_matchingBytes_2400(matchingBytes[2400]),
.io_matchingBytes_2401(matchingBytes[2401]),
.io_matchingBytes_2402(matchingBytes[2402]),
.io_matchingBytes_2403(matchingBytes[2403]),
.io_matchingBytes_2404(matchingBytes[2404]),
.io_matchingBytes_2405(matchingBytes[2405]),
.io_matchingBytes_2406(matchingBytes[2406]),
.io_matchingBytes_2407(matchingBytes[2407]),
.io_matchingBytes_2408(matchingBytes[2408]),
.io_matchingBytes_2409(matchingBytes[2409]),
.io_matchingBytes_2410(matchingBytes[2410]),
.io_matchingBytes_2411(matchingBytes[2411]),
.io_matchingBytes_2412(matchingBytes[2412]),
.io_matchingBytes_2413(matchingBytes[2413]),
.io_matchingBytes_2414(matchingBytes[2414]),
.io_matchingBytes_2415(matchingBytes[2415]),
.io_matchingBytes_2416(matchingBytes[2416]),
.io_matchingBytes_2417(matchingBytes[2417]),
.io_matchingBytes_2418(matchingBytes[2418]),
.io_matchingBytes_2419(matchingBytes[2419]),
.io_matchingBytes_2420(matchingBytes[2420]),
.io_matchingBytes_2421(matchingBytes[2421]),
.io_matchingBytes_2422(matchingBytes[2422]),
.io_matchingBytes_2423(matchingBytes[2423]),
.io_matchingBytes_2424(matchingBytes[2424]),
.io_matchingBytes_2425(matchingBytes[2425]),
.io_matchingBytes_2426(matchingBytes[2426]),
.io_matchingBytes_2427(matchingBytes[2427]),
.io_matchingBytes_2428(matchingBytes[2428]),
.io_matchingBytes_2429(matchingBytes[2429]),
.io_matchingBytes_2430(matchingBytes[2430]),
.io_matchingBytes_2431(matchingBytes[2431]),
.io_matchingBytes_2432(matchingBytes[2432]),
.io_matchingBytes_2433(matchingBytes[2433]),
.io_matchingBytes_2434(matchingBytes[2434]),
.io_matchingBytes_2435(matchingBytes[2435]),
.io_matchingBytes_2436(matchingBytes[2436]),
.io_matchingBytes_2437(matchingBytes[2437]),
.io_matchingBytes_2438(matchingBytes[2438]),
.io_matchingBytes_2439(matchingBytes[2439]),
.io_matchingBytes_2440(matchingBytes[2440]),
.io_matchingBytes_2441(matchingBytes[2441]),
.io_matchingBytes_2442(matchingBytes[2442]),
.io_matchingBytes_2443(matchingBytes[2443]),
.io_matchingBytes_2444(matchingBytes[2444]),
.io_matchingBytes_2445(matchingBytes[2445]),
.io_matchingBytes_2446(matchingBytes[2446]),
.io_matchingBytes_2447(matchingBytes[2447]),
.io_matchingBytes_2448(matchingBytes[2448]),
.io_matchingBytes_2449(matchingBytes[2449]),
.io_matchingBytes_2450(matchingBytes[2450]),
.io_matchingBytes_2451(matchingBytes[2451]),
.io_matchingBytes_2452(matchingBytes[2452]),
.io_matchingBytes_2453(matchingBytes[2453]),
.io_matchingBytes_2454(matchingBytes[2454]),
.io_matchingBytes_2455(matchingBytes[2455]),
.io_matchingBytes_2456(matchingBytes[2456]),
.io_matchingBytes_2457(matchingBytes[2457]),
.io_matchingBytes_2458(matchingBytes[2458]),
.io_matchingBytes_2459(matchingBytes[2459]),
.io_matchingBytes_2460(matchingBytes[2460]),
.io_matchingBytes_2461(matchingBytes[2461]),
.io_matchingBytes_2462(matchingBytes[2462]),
.io_matchingBytes_2463(matchingBytes[2463]),
.io_matchingBytes_2464(matchingBytes[2464]),
.io_matchingBytes_2465(matchingBytes[2465]),
.io_matchingBytes_2466(matchingBytes[2466]),
.io_matchingBytes_2467(matchingBytes[2467]),
.io_matchingBytes_2468(matchingBytes[2468]),
.io_matchingBytes_2469(matchingBytes[2469]),
.io_matchingBytes_2470(matchingBytes[2470]),
.io_matchingBytes_2471(matchingBytes[2471]),
.io_matchingBytes_2472(matchingBytes[2472]),
.io_matchingBytes_2473(matchingBytes[2473]),
.io_matchingBytes_2474(matchingBytes[2474]),
.io_matchingBytes_2475(matchingBytes[2475]),
.io_matchingBytes_2476(matchingBytes[2476]),
.io_matchingBytes_2477(matchingBytes[2477]),
.io_matchingBytes_2478(matchingBytes[2478]),
.io_matchingBytes_2479(matchingBytes[2479]),
.io_matchingBytes_2480(matchingBytes[2480]),
.io_matchingBytes_2481(matchingBytes[2481]),
.io_matchingBytes_2482(matchingBytes[2482]),
.io_matchingBytes_2483(matchingBytes[2483]),
.io_matchingBytes_2484(matchingBytes[2484]),
.io_matchingBytes_2485(matchingBytes[2485]),
.io_matchingBytes_2486(matchingBytes[2486]),
.io_matchingBytes_2487(matchingBytes[2487]),
.io_matchingBytes_2488(matchingBytes[2488]),
.io_matchingBytes_2489(matchingBytes[2489]),
.io_matchingBytes_2490(matchingBytes[2490]),
.io_matchingBytes_2491(matchingBytes[2491]),
.io_matchingBytes_2492(matchingBytes[2492]),
.io_matchingBytes_2493(matchingBytes[2493]),
.io_matchingBytes_2494(matchingBytes[2494]),
.io_matchingBytes_2495(matchingBytes[2495]),
.io_matchingBytes_2496(matchingBytes[2496]),
.io_matchingBytes_2497(matchingBytes[2497]),
.io_matchingBytes_2498(matchingBytes[2498]),
.io_matchingBytes_2499(matchingBytes[2499]),
.io_matchingBytes_2500(matchingBytes[2500]),
.io_matchingBytes_2501(matchingBytes[2501]),
.io_matchingBytes_2502(matchingBytes[2502]),
.io_matchingBytes_2503(matchingBytes[2503]),
.io_matchingBytes_2504(matchingBytes[2504]),
.io_matchingBytes_2505(matchingBytes[2505]),
.io_matchingBytes_2506(matchingBytes[2506]),
.io_matchingBytes_2507(matchingBytes[2507]),
.io_matchingBytes_2508(matchingBytes[2508]),
.io_matchingBytes_2509(matchingBytes[2509]),
.io_matchingBytes_2510(matchingBytes[2510]),
.io_matchingBytes_2511(matchingBytes[2511]),
.io_matchingBytes_2512(matchingBytes[2512]),
.io_matchingBytes_2513(matchingBytes[2513]),
.io_matchingBytes_2514(matchingBytes[2514]),
.io_matchingBytes_2515(matchingBytes[2515]),
.io_matchingBytes_2516(matchingBytes[2516]),
.io_matchingBytes_2517(matchingBytes[2517]),
.io_matchingBytes_2518(matchingBytes[2518]),
.io_matchingBytes_2519(matchingBytes[2519]),
.io_matchingBytes_2520(matchingBytes[2520]),
.io_matchingBytes_2521(matchingBytes[2521]),
.io_matchingBytes_2522(matchingBytes[2522]),
.io_matchingBytes_2523(matchingBytes[2523]),
.io_matchingBytes_2524(matchingBytes[2524]),
.io_matchingBytes_2525(matchingBytes[2525]),
.io_matchingBytes_2526(matchingBytes[2526]),
.io_matchingBytes_2527(matchingBytes[2527]),
.io_matchingBytes_2528(matchingBytes[2528]),
.io_matchingBytes_2529(matchingBytes[2529]),
.io_matchingBytes_2530(matchingBytes[2530]),
.io_matchingBytes_2531(matchingBytes[2531]),
.io_matchingBytes_2532(matchingBytes[2532]),
.io_matchingBytes_2533(matchingBytes[2533]),
.io_matchingBytes_2534(matchingBytes[2534]),
.io_matchingBytes_2535(matchingBytes[2535]),
.io_matchingBytes_2536(matchingBytes[2536]),
.io_matchingBytes_2537(matchingBytes[2537]),
.io_matchingBytes_2538(matchingBytes[2538]),
.io_matchingBytes_2539(matchingBytes[2539]),
.io_matchingBytes_2540(matchingBytes[2540]),
.io_matchingBytes_2541(matchingBytes[2541]),
.io_matchingBytes_2542(matchingBytes[2542]),
.io_matchingBytes_2543(matchingBytes[2543]),
.io_matchingBytes_2544(matchingBytes[2544]),
.io_matchingBytes_2545(matchingBytes[2545]),
.io_matchingBytes_2546(matchingBytes[2546]),
.io_matchingBytes_2547(matchingBytes[2547]),
.io_matchingBytes_2548(matchingBytes[2548]),
.io_matchingBytes_2549(matchingBytes[2549]),
.io_matchingBytes_2550(matchingBytes[2550]),
.io_matchingBytes_2551(matchingBytes[2551]),
.io_matchingBytes_2552(matchingBytes[2552]),
.io_matchingBytes_2553(matchingBytes[2553]),
.io_matchingBytes_2554(matchingBytes[2554]),
.io_matchingBytes_2555(matchingBytes[2555]),
.io_matchingBytes_2556(matchingBytes[2556]),
.io_matchingBytes_2557(matchingBytes[2557]),
.io_matchingBytes_2558(matchingBytes[2558]),
.io_matchingBytes_2559(matchingBytes[2559]),
.io_matchingBytes_2560(matchingBytes[2560]),
.io_matchingBytes_2561(matchingBytes[2561]),
.io_matchingBytes_2562(matchingBytes[2562]),
.io_matchingBytes_2563(matchingBytes[2563]),
.io_matchingBytes_2564(matchingBytes[2564]),
.io_matchingBytes_2565(matchingBytes[2565]),
.io_matchingBytes_2566(matchingBytes[2566]),
.io_matchingBytes_2567(matchingBytes[2567]),
.io_matchingBytes_2568(matchingBytes[2568]),
.io_matchingBytes_2569(matchingBytes[2569]),
.io_matchingBytes_2570(matchingBytes[2570]),
.io_matchingBytes_2571(matchingBytes[2571]),
.io_matchingBytes_2572(matchingBytes[2572]),
.io_matchingBytes_2573(matchingBytes[2573]),
.io_matchingBytes_2574(matchingBytes[2574]),
.io_matchingBytes_2575(matchingBytes[2575]),
.io_matchingBytes_2576(matchingBytes[2576]),
.io_matchingBytes_2577(matchingBytes[2577]),
.io_matchingBytes_2578(matchingBytes[2578]),
.io_matchingBytes_2579(matchingBytes[2579]),
.io_matchingBytes_2580(matchingBytes[2580]),
.io_matchingBytes_2581(matchingBytes[2581]),
.io_matchingBytes_2582(matchingBytes[2582]),
.io_matchingBytes_2583(matchingBytes[2583]),
.io_matchingBytes_2584(matchingBytes[2584]),
.io_matchingBytes_2585(matchingBytes[2585]),
.io_matchingBytes_2586(matchingBytes[2586]),
.io_matchingBytes_2587(matchingBytes[2587]),
.io_matchingBytes_2588(matchingBytes[2588]),
.io_matchingBytes_2589(matchingBytes[2589]),
.io_matchingBytes_2590(matchingBytes[2590]),
.io_matchingBytes_2591(matchingBytes[2591]),
.io_matchingBytes_2592(matchingBytes[2592]),
.io_matchingBytes_2593(matchingBytes[2593]),
.io_matchingBytes_2594(matchingBytes[2594]),
.io_matchingBytes_2595(matchingBytes[2595]),
.io_matchingBytes_2596(matchingBytes[2596]),
.io_matchingBytes_2597(matchingBytes[2597]),
.io_matchingBytes_2598(matchingBytes[2598]),
.io_matchingBytes_2599(matchingBytes[2599]),
.io_matchingBytes_2600(matchingBytes[2600]),
.io_matchingBytes_2601(matchingBytes[2601]),
.io_matchingBytes_2602(matchingBytes[2602]),
.io_matchingBytes_2603(matchingBytes[2603]),
.io_matchingBytes_2604(matchingBytes[2604]),
.io_matchingBytes_2605(matchingBytes[2605]),
.io_matchingBytes_2606(matchingBytes[2606]),
.io_matchingBytes_2607(matchingBytes[2607]),
.io_matchingBytes_2608(matchingBytes[2608]),
.io_matchingBytes_2609(matchingBytes[2609]),
.io_matchingBytes_2610(matchingBytes[2610]),
.io_matchingBytes_2611(matchingBytes[2611]),
.io_matchingBytes_2612(matchingBytes[2612]),
.io_matchingBytes_2613(matchingBytes[2613]),
.io_matchingBytes_2614(matchingBytes[2614]),
.io_matchingBytes_2615(matchingBytes[2615]),
.io_matchingBytes_2616(matchingBytes[2616]),
.io_matchingBytes_2617(matchingBytes[2617]),
.io_matchingBytes_2618(matchingBytes[2618]),
.io_matchingBytes_2619(matchingBytes[2619]),
.io_matchingBytes_2620(matchingBytes[2620]),
.io_matchingBytes_2621(matchingBytes[2621]),
.io_matchingBytes_2622(matchingBytes[2622]),
.io_matchingBytes_2623(matchingBytes[2623]),
.io_matchingBytes_2624(matchingBytes[2624]),
.io_matchingBytes_2625(matchingBytes[2625]),
.io_matchingBytes_2626(matchingBytes[2626]),
.io_matchingBytes_2627(matchingBytes[2627]),
.io_matchingBytes_2628(matchingBytes[2628]),
.io_matchingBytes_2629(matchingBytes[2629]),
.io_matchingBytes_2630(matchingBytes[2630]),
.io_matchingBytes_2631(matchingBytes[2631]),
.io_matchingBytes_2632(matchingBytes[2632]),
.io_matchingBytes_2633(matchingBytes[2633]),
.io_matchingBytes_2634(matchingBytes[2634]),
.io_matchingBytes_2635(matchingBytes[2635]),
.io_matchingBytes_2636(matchingBytes[2636]),
.io_matchingBytes_2637(matchingBytes[2637]),
.io_matchingBytes_2638(matchingBytes[2638]),
.io_matchingBytes_2639(matchingBytes[2639]),
.io_matchingBytes_2640(matchingBytes[2640]),
.io_matchingBytes_2641(matchingBytes[2641]),
.io_matchingBytes_2642(matchingBytes[2642]),
.io_matchingBytes_2643(matchingBytes[2643]),
.io_matchingBytes_2644(matchingBytes[2644]),
.io_matchingBytes_2645(matchingBytes[2645]),
.io_matchingBytes_2646(matchingBytes[2646]),
.io_matchingBytes_2647(matchingBytes[2647]),
.io_matchingBytes_2648(matchingBytes[2648]),
.io_matchingBytes_2649(matchingBytes[2649]),
.io_matchingBytes_2650(matchingBytes[2650]),
.io_matchingBytes_2651(matchingBytes[2651]),
.io_matchingBytes_2652(matchingBytes[2652]),
.io_matchingBytes_2653(matchingBytes[2653]),
.io_matchingBytes_2654(matchingBytes[2654]),
.io_matchingBytes_2655(matchingBytes[2655]),
.io_matchingBytes_2656(matchingBytes[2656]),
.io_matchingBytes_2657(matchingBytes[2657]),
.io_matchingBytes_2658(matchingBytes[2658]),
.io_matchingBytes_2659(matchingBytes[2659]),
.io_matchingBytes_2660(matchingBytes[2660]),
.io_matchingBytes_2661(matchingBytes[2661]),
.io_matchingBytes_2662(matchingBytes[2662]),
.io_matchingBytes_2663(matchingBytes[2663]),
.io_matchingBytes_2664(matchingBytes[2664]),
.io_matchingBytes_2665(matchingBytes[2665]),
.io_matchingBytes_2666(matchingBytes[2666]),
.io_matchingBytes_2667(matchingBytes[2667]),
.io_matchingBytes_2668(matchingBytes[2668]),
.io_matchingBytes_2669(matchingBytes[2669]),
.io_matchingBytes_2670(matchingBytes[2670]),
.io_matchingBytes_2671(matchingBytes[2671]),
.io_matchingBytes_2672(matchingBytes[2672]),
.io_matchingBytes_2673(matchingBytes[2673]),
.io_matchingBytes_2674(matchingBytes[2674]),
.io_matchingBytes_2675(matchingBytes[2675]),
.io_matchingBytes_2676(matchingBytes[2676]),
.io_matchingBytes_2677(matchingBytes[2677]),
.io_matchingBytes_2678(matchingBytes[2678]),
.io_matchingBytes_2679(matchingBytes[2679]),
.io_matchingBytes_2680(matchingBytes[2680]),
.io_matchingBytes_2681(matchingBytes[2681]),
.io_matchingBytes_2682(matchingBytes[2682]),
.io_matchingBytes_2683(matchingBytes[2683]),
.io_matchingBytes_2684(matchingBytes[2684]),
.io_matchingBytes_2685(matchingBytes[2685]),
.io_matchingBytes_2686(matchingBytes[2686]),
.io_matchingBytes_2687(matchingBytes[2687]),
.io_matchingBytes_2688(matchingBytes[2688]),
.io_matchingBytes_2689(matchingBytes[2689]),
.io_matchingBytes_2690(matchingBytes[2690]),
.io_matchingBytes_2691(matchingBytes[2691]),
.io_matchingBytes_2692(matchingBytes[2692]),
.io_matchingBytes_2693(matchingBytes[2693]),
.io_matchingBytes_2694(matchingBytes[2694]),
.io_matchingBytes_2695(matchingBytes[2695]),
.io_matchingBytes_2696(matchingBytes[2696]),
.io_matchingBytes_2697(matchingBytes[2697]),
.io_matchingBytes_2698(matchingBytes[2698]),
.io_matchingBytes_2699(matchingBytes[2699]),
.io_matchingBytes_2700(matchingBytes[2700]),
.io_matchingBytes_2701(matchingBytes[2701]),
.io_matchingBytes_2702(matchingBytes[2702]),
.io_matchingBytes_2703(matchingBytes[2703]),
.io_matchingBytes_2704(matchingBytes[2704]),
.io_matchingBytes_2705(matchingBytes[2705]),
.io_matchingBytes_2706(matchingBytes[2706]),
.io_matchingBytes_2707(matchingBytes[2707]),
.io_matchingBytes_2708(matchingBytes[2708]),
.io_matchingBytes_2709(matchingBytes[2709]),
.io_matchingBytes_2710(matchingBytes[2710]),
.io_matchingBytes_2711(matchingBytes[2711]),
.io_matchingBytes_2712(matchingBytes[2712]),
.io_matchingBytes_2713(matchingBytes[2713]),
.io_matchingBytes_2714(matchingBytes[2714]),
.io_matchingBytes_2715(matchingBytes[2715]),
.io_matchingBytes_2716(matchingBytes[2716]),
.io_matchingBytes_2717(matchingBytes[2717]),
.io_matchingBytes_2718(matchingBytes[2718]),
.io_matchingBytes_2719(matchingBytes[2719]),
.io_matchingBytes_2720(matchingBytes[2720]),
.io_matchingBytes_2721(matchingBytes[2721]),
.io_matchingBytes_2722(matchingBytes[2722]),
.io_matchingBytes_2723(matchingBytes[2723]),
.io_matchingBytes_2724(matchingBytes[2724]),
.io_matchingBytes_2725(matchingBytes[2725]),
.io_matchingBytes_2726(matchingBytes[2726]),
.io_matchingBytes_2727(matchingBytes[2727]),
.io_matchingBytes_2728(matchingBytes[2728]),
.io_matchingBytes_2729(matchingBytes[2729]),
.io_matchingBytes_2730(matchingBytes[2730]),
.io_matchingBytes_2731(matchingBytes[2731]),
.io_matchingBytes_2732(matchingBytes[2732]),
.io_matchingBytes_2733(matchingBytes[2733]),
.io_matchingBytes_2734(matchingBytes[2734]),
.io_matchingBytes_2735(matchingBytes[2735]),
.io_matchingBytes_2736(matchingBytes[2736]),
.io_matchingBytes_2737(matchingBytes[2737]),
.io_matchingBytes_2738(matchingBytes[2738]),
.io_matchingBytes_2739(matchingBytes[2739]),
.io_matchingBytes_2740(matchingBytes[2740]),
.io_matchingBytes_2741(matchingBytes[2741]),
.io_matchingBytes_2742(matchingBytes[2742]),
.io_matchingBytes_2743(matchingBytes[2743]),
.io_matchingBytes_2744(matchingBytes[2744]),
.io_matchingBytes_2745(matchingBytes[2745]),
.io_matchingBytes_2746(matchingBytes[2746]),
.io_matchingBytes_2747(matchingBytes[2747]),
.io_matchingBytes_2748(matchingBytes[2748]),
.io_matchingBytes_2749(matchingBytes[2749]),
.io_matchingBytes_2750(matchingBytes[2750]),
.io_matchingBytes_2751(matchingBytes[2751]),
.io_matchingBytes_2752(matchingBytes[2752]),
.io_matchingBytes_2753(matchingBytes[2753]),
.io_matchingBytes_2754(matchingBytes[2754]),
.io_matchingBytes_2755(matchingBytes[2755]),
.io_matchingBytes_2756(matchingBytes[2756]),
.io_matchingBytes_2757(matchingBytes[2757]),
.io_matchingBytes_2758(matchingBytes[2758]),
.io_matchingBytes_2759(matchingBytes[2759]),
.io_matchingBytes_2760(matchingBytes[2760]),
.io_matchingBytes_2761(matchingBytes[2761]),
.io_matchingBytes_2762(matchingBytes[2762]),
.io_matchingBytes_2763(matchingBytes[2763]),
.io_matchingBytes_2764(matchingBytes[2764]),
.io_matchingBytes_2765(matchingBytes[2765]),
.io_matchingBytes_2766(matchingBytes[2766]),
.io_matchingBytes_2767(matchingBytes[2767]),
.io_matchingBytes_2768(matchingBytes[2768]),
.io_matchingBytes_2769(matchingBytes[2769]),
.io_matchingBytes_2770(matchingBytes[2770]),
.io_matchingBytes_2771(matchingBytes[2771]),
.io_matchingBytes_2772(matchingBytes[2772]),
.io_matchingBytes_2773(matchingBytes[2773]),
.io_matchingBytes_2774(matchingBytes[2774]),
.io_matchingBytes_2775(matchingBytes[2775]),
.io_matchingBytes_2776(matchingBytes[2776]),
.io_matchingBytes_2777(matchingBytes[2777]),
.io_matchingBytes_2778(matchingBytes[2778]),
.io_matchingBytes_2779(matchingBytes[2779]),
.io_matchingBytes_2780(matchingBytes[2780]),
.io_matchingBytes_2781(matchingBytes[2781]),
.io_matchingBytes_2782(matchingBytes[2782]),
.io_matchingBytes_2783(matchingBytes[2783]),
.io_matchingBytes_2784(matchingBytes[2784]),
.io_matchingBytes_2785(matchingBytes[2785]),
.io_matchingBytes_2786(matchingBytes[2786]),
.io_matchingBytes_2787(matchingBytes[2787]),
.io_matchingBytes_2788(matchingBytes[2788]),
.io_matchingBytes_2789(matchingBytes[2789]),
.io_matchingBytes_2790(matchingBytes[2790]),
.io_matchingBytes_2791(matchingBytes[2791]),
.io_matchingBytes_2792(matchingBytes[2792]),
.io_matchingBytes_2793(matchingBytes[2793]),
.io_matchingBytes_2794(matchingBytes[2794]),
.io_matchingBytes_2795(matchingBytes[2795]),
.io_matchingBytes_2796(matchingBytes[2796]),
.io_matchingBytes_2797(matchingBytes[2797]),
.io_matchingBytes_2798(matchingBytes[2798]),
.io_matchingBytes_2799(matchingBytes[2799]),
.io_matchingBytes_2800(matchingBytes[2800]),
.io_matchingBytes_2801(matchingBytes[2801]),
.io_matchingBytes_2802(matchingBytes[2802]),
.io_matchingBytes_2803(matchingBytes[2803]),
.io_matchingBytes_2804(matchingBytes[2804]),
.io_matchingBytes_2805(matchingBytes[2805]),
.io_matchingBytes_2806(matchingBytes[2806]),
.io_matchingBytes_2807(matchingBytes[2807]),
.io_matchingBytes_2808(matchingBytes[2808]),
.io_matchingBytes_2809(matchingBytes[2809]),
.io_matchingBytes_2810(matchingBytes[2810]),
.io_matchingBytes_2811(matchingBytes[2811]),
.io_matchingBytes_2812(matchingBytes[2812]),
.io_matchingBytes_2813(matchingBytes[2813]),
.io_matchingBytes_2814(matchingBytes[2814]),
.io_matchingBytes_2815(matchingBytes[2815]),
.io_matchingBytes_2816(matchingBytes[2816]),
.io_matchingBytes_2817(matchingBytes[2817]),
.io_matchingBytes_2818(matchingBytes[2818]),
.io_matchingBytes_2819(matchingBytes[2819]),
.io_matchingBytes_2820(matchingBytes[2820]),
.io_matchingBytes_2821(matchingBytes[2821]),
.io_matchingBytes_2822(matchingBytes[2822]),
.io_matchingBytes_2823(matchingBytes[2823]),
.io_matchingBytes_2824(matchingBytes[2824]),
.io_matchingBytes_2825(matchingBytes[2825]),
.io_matchingBytes_2826(matchingBytes[2826]),
.io_matchingBytes_2827(matchingBytes[2827]),
.io_matchingBytes_2828(matchingBytes[2828]),
.io_matchingBytes_2829(matchingBytes[2829]),
.io_matchingBytes_2830(matchingBytes[2830]),
.io_matchingBytes_2831(matchingBytes[2831]),
.io_matchingBytes_2832(matchingBytes[2832]),
.io_matchingBytes_2833(matchingBytes[2833]),
.io_matchingBytes_2834(matchingBytes[2834]),
.io_matchingBytes_2835(matchingBytes[2835]),
.io_matchingBytes_2836(matchingBytes[2836]),
.io_matchingBytes_2837(matchingBytes[2837]),
.io_matchingBytes_2838(matchingBytes[2838]),
.io_matchingBytes_2839(matchingBytes[2839]),
.io_matchingBytes_2840(matchingBytes[2840]),
.io_matchingBytes_2841(matchingBytes[2841]),
.io_matchingBytes_2842(matchingBytes[2842]),
.io_matchingBytes_2843(matchingBytes[2843]),
.io_matchingBytes_2844(matchingBytes[2844]),
.io_matchingBytes_2845(matchingBytes[2845]),
.io_matchingBytes_2846(matchingBytes[2846]),
.io_matchingBytes_2847(matchingBytes[2847]),
.io_matchingBytes_2848(matchingBytes[2848]),
.io_matchingBytes_2849(matchingBytes[2849]),
.io_matchingBytes_2850(matchingBytes[2850]),
.io_matchingBytes_2851(matchingBytes[2851]),
.io_matchingBytes_2852(matchingBytes[2852]),
.io_matchingBytes_2853(matchingBytes[2853]),
.io_matchingBytes_2854(matchingBytes[2854]),
.io_matchingBytes_2855(matchingBytes[2855]),
.io_matchingBytes_2856(matchingBytes[2856]),
.io_matchingBytes_2857(matchingBytes[2857]),
.io_matchingBytes_2858(matchingBytes[2858]),
.io_matchingBytes_2859(matchingBytes[2859]),
.io_matchingBytes_2860(matchingBytes[2860]),
.io_matchingBytes_2861(matchingBytes[2861]),
.io_matchingBytes_2862(matchingBytes[2862]),
.io_matchingBytes_2863(matchingBytes[2863]),
.io_matchingBytes_2864(matchingBytes[2864]),
.io_matchingBytes_2865(matchingBytes[2865]),
.io_matchingBytes_2866(matchingBytes[2866]),
.io_matchingBytes_2867(matchingBytes[2867]),
.io_matchingBytes_2868(matchingBytes[2868]),
.io_matchingBytes_2869(matchingBytes[2869]),
.io_matchingBytes_2870(matchingBytes[2870]),
.io_matchingBytes_2871(matchingBytes[2871]),
.io_matchingBytes_2872(matchingBytes[2872]),
.io_matchingBytes_2873(matchingBytes[2873]),
.io_matchingBytes_2874(matchingBytes[2874]),
.io_matchingBytes_2875(matchingBytes[2875]),
.io_matchingBytes_2876(matchingBytes[2876]),
.io_matchingBytes_2877(matchingBytes[2877]),
.io_matchingBytes_2878(matchingBytes[2878]),
.io_matchingBytes_2879(matchingBytes[2879]),
.io_matchingBytes_2880(matchingBytes[2880]),
.io_matchingBytes_2881(matchingBytes[2881]),
.io_matchingBytes_2882(matchingBytes[2882]),
.io_matchingBytes_2883(matchingBytes[2883]),
.io_matchingBytes_2884(matchingBytes[2884]),
.io_matchingBytes_2885(matchingBytes[2885]),
.io_matchingBytes_2886(matchingBytes[2886]),
.io_matchingBytes_2887(matchingBytes[2887]),
.io_matchingBytes_2888(matchingBytes[2888]),
.io_matchingBytes_2889(matchingBytes[2889]),
.io_matchingBytes_2890(matchingBytes[2890]),
.io_matchingBytes_2891(matchingBytes[2891]),
.io_matchingBytes_2892(matchingBytes[2892]),
.io_matchingBytes_2893(matchingBytes[2893]),
.io_matchingBytes_2894(matchingBytes[2894]),
.io_matchingBytes_2895(matchingBytes[2895]),
.io_matchingBytes_2896(matchingBytes[2896]),
.io_matchingBytes_2897(matchingBytes[2897]),
.io_matchingBytes_2898(matchingBytes[2898]),
.io_matchingBytes_2899(matchingBytes[2899]),
.io_matchingBytes_2900(matchingBytes[2900]),
.io_matchingBytes_2901(matchingBytes[2901]),
.io_matchingBytes_2902(matchingBytes[2902]),
.io_matchingBytes_2903(matchingBytes[2903]),
.io_matchingBytes_2904(matchingBytes[2904]),
.io_matchingBytes_2905(matchingBytes[2905]),
.io_matchingBytes_2906(matchingBytes[2906]),
.io_matchingBytes_2907(matchingBytes[2907]),
.io_matchingBytes_2908(matchingBytes[2908]),
.io_matchingBytes_2909(matchingBytes[2909]),
.io_matchingBytes_2910(matchingBytes[2910]),
.io_matchingBytes_2911(matchingBytes[2911]),
.io_matchingBytes_2912(matchingBytes[2912]),
.io_matchingBytes_2913(matchingBytes[2913]),
.io_matchingBytes_2914(matchingBytes[2914]),
.io_matchingBytes_2915(matchingBytes[2915]),
.io_matchingBytes_2916(matchingBytes[2916]),
.io_matchingBytes_2917(matchingBytes[2917]),
.io_matchingBytes_2918(matchingBytes[2918]),
.io_matchingBytes_2919(matchingBytes[2919]),
.io_matchingBytes_2920(matchingBytes[2920]),
.io_matchingBytes_2921(matchingBytes[2921]),
.io_matchingBytes_2922(matchingBytes[2922]),
.io_matchingBytes_2923(matchingBytes[2923]),
.io_matchingBytes_2924(matchingBytes[2924]),
.io_matchingBytes_2925(matchingBytes[2925]),
.io_matchingBytes_2926(matchingBytes[2926]),
.io_matchingBytes_2927(matchingBytes[2927]),
.io_matchingBytes_2928(matchingBytes[2928]),
.io_matchingBytes_2929(matchingBytes[2929]),
.io_matchingBytes_2930(matchingBytes[2930]),
.io_matchingBytes_2931(matchingBytes[2931]),
.io_matchingBytes_2932(matchingBytes[2932]),
.io_matchingBytes_2933(matchingBytes[2933]),
.io_matchingBytes_2934(matchingBytes[2934]),
.io_matchingBytes_2935(matchingBytes[2935]),
.io_matchingBytes_2936(matchingBytes[2936]),
.io_matchingBytes_2937(matchingBytes[2937]),
.io_matchingBytes_2938(matchingBytes[2938]),
.io_matchingBytes_2939(matchingBytes[2939]),
.io_matchingBytes_2940(matchingBytes[2940]),
.io_matchingBytes_2941(matchingBytes[2941]),
.io_matchingBytes_2942(matchingBytes[2942]),
.io_matchingBytes_2943(matchingBytes[2943]),
.io_matchingBytes_2944(matchingBytes[2944]),
.io_matchingBytes_2945(matchingBytes[2945]),
.io_matchingBytes_2946(matchingBytes[2946]),
.io_matchingBytes_2947(matchingBytes[2947]),
.io_matchingBytes_2948(matchingBytes[2948]),
.io_matchingBytes_2949(matchingBytes[2949]),
.io_matchingBytes_2950(matchingBytes[2950]),
.io_matchingBytes_2951(matchingBytes[2951]),
.io_matchingBytes_2952(matchingBytes[2952]),
.io_matchingBytes_2953(matchingBytes[2953]),
.io_matchingBytes_2954(matchingBytes[2954]),
.io_matchingBytes_2955(matchingBytes[2955]),
.io_matchingBytes_2956(matchingBytes[2956]),
.io_matchingBytes_2957(matchingBytes[2957]),
.io_matchingBytes_2958(matchingBytes[2958]),
.io_matchingBytes_2959(matchingBytes[2959]),
.io_matchingBytes_2960(matchingBytes[2960]),
.io_matchingBytes_2961(matchingBytes[2961]),
.io_matchingBytes_2962(matchingBytes[2962]),
.io_matchingBytes_2963(matchingBytes[2963]),
.io_matchingBytes_2964(matchingBytes[2964]),
.io_matchingBytes_2965(matchingBytes[2965]),
.io_matchingBytes_2966(matchingBytes[2966]),
.io_matchingBytes_2967(matchingBytes[2967]),
.io_matchingBytes_2968(matchingBytes[2968]),
.io_matchingBytes_2969(matchingBytes[2969]),
.io_matchingBytes_2970(matchingBytes[2970]),
.io_matchingBytes_2971(matchingBytes[2971]),
.io_matchingBytes_2972(matchingBytes[2972]),
.io_matchingBytes_2973(matchingBytes[2973]),
.io_matchingBytes_2974(matchingBytes[2974]),
.io_matchingBytes_2975(matchingBytes[2975]),
.io_matchingBytes_2976(matchingBytes[2976]),
.io_matchingBytes_2977(matchingBytes[2977]),
.io_matchingBytes_2978(matchingBytes[2978]),
.io_matchingBytes_2979(matchingBytes[2979]),
.io_matchingBytes_2980(matchingBytes[2980]),
.io_matchingBytes_2981(matchingBytes[2981]),
.io_matchingBytes_2982(matchingBytes[2982]),
.io_matchingBytes_2983(matchingBytes[2983]),
.io_matchingBytes_2984(matchingBytes[2984]),
.io_matchingBytes_2985(matchingBytes[2985]),
.io_matchingBytes_2986(matchingBytes[2986]),
.io_matchingBytes_2987(matchingBytes[2987]),
.io_matchingBytes_2988(matchingBytes[2988]),
.io_matchingBytes_2989(matchingBytes[2989]),
.io_matchingBytes_2990(matchingBytes[2990]),
.io_matchingBytes_2991(matchingBytes[2991]),
.io_matchingBytes_2992(matchingBytes[2992]),
.io_matchingBytes_2993(matchingBytes[2993]),
.io_matchingBytes_2994(matchingBytes[2994]),
.io_matchingBytes_2995(matchingBytes[2995]),
.io_matchingBytes_2996(matchingBytes[2996]),
.io_matchingBytes_2997(matchingBytes[2997]),
.io_matchingBytes_2998(matchingBytes[2998]),
.io_matchingBytes_2999(matchingBytes[2999]),
.io_matchingBytes_3000(matchingBytes[3000]),
.io_matchingBytes_3001(matchingBytes[3001]),
.io_matchingBytes_3002(matchingBytes[3002]),
.io_matchingBytes_3003(matchingBytes[3003]),
.io_matchingBytes_3004(matchingBytes[3004]),
.io_matchingBytes_3005(matchingBytes[3005]),
.io_matchingBytes_3006(matchingBytes[3006]),
.io_matchingBytes_3007(matchingBytes[3007]),
.io_matchingBytes_3008(matchingBytes[3008]),
.io_matchingBytes_3009(matchingBytes[3009]),
.io_matchingBytes_3010(matchingBytes[3010]),
.io_matchingBytes_3011(matchingBytes[3011]),
.io_matchingBytes_3012(matchingBytes[3012]),
.io_matchingBytes_3013(matchingBytes[3013]),
.io_matchingBytes_3014(matchingBytes[3014]),
.io_matchingBytes_3015(matchingBytes[3015]),
.io_matchingBytes_3016(matchingBytes[3016]),
.io_matchingBytes_3017(matchingBytes[3017]),
.io_matchingBytes_3018(matchingBytes[3018]),
.io_matchingBytes_3019(matchingBytes[3019]),
.io_matchingBytes_3020(matchingBytes[3020]),
.io_matchingBytes_3021(matchingBytes[3021]),
.io_matchingBytes_3022(matchingBytes[3022]),
.io_matchingBytes_3023(matchingBytes[3023]),
.io_matchingBytes_3024(matchingBytes[3024]),
.io_matchingBytes_3025(matchingBytes[3025]),
.io_matchingBytes_3026(matchingBytes[3026]),
.io_matchingBytes_3027(matchingBytes[3027]),
.io_matchingBytes_3028(matchingBytes[3028]),
.io_matchingBytes_3029(matchingBytes[3029]),
.io_matchingBytes_3030(matchingBytes[3030]),
.io_matchingBytes_3031(matchingBytes[3031]),
.io_matchingBytes_3032(matchingBytes[3032]),
.io_matchingBytes_3033(matchingBytes[3033]),
.io_matchingBytes_3034(matchingBytes[3034]),
.io_matchingBytes_3035(matchingBytes[3035]),
.io_matchingBytes_3036(matchingBytes[3036]),
.io_matchingBytes_3037(matchingBytes[3037]),
.io_matchingBytes_3038(matchingBytes[3038]),
.io_matchingBytes_3039(matchingBytes[3039]),
.io_matchingBytes_3040(matchingBytes[3040]),
.io_matchingBytes_3041(matchingBytes[3041]),
.io_matchingBytes_3042(matchingBytes[3042]),
.io_matchingBytes_3043(matchingBytes[3043]),
.io_matchingBytes_3044(matchingBytes[3044]),
.io_matchingBytes_3045(matchingBytes[3045]),
.io_matchingBytes_3046(matchingBytes[3046]),
.io_matchingBytes_3047(matchingBytes[3047]),
.io_matchingBytes_3048(matchingBytes[3048]),
.io_matchingBytes_3049(matchingBytes[3049]),
.io_matchingBytes_3050(matchingBytes[3050]),
.io_matchingBytes_3051(matchingBytes[3051]),
.io_matchingBytes_3052(matchingBytes[3052]),
.io_matchingBytes_3053(matchingBytes[3053]),
.io_matchingBytes_3054(matchingBytes[3054]),
.io_matchingBytes_3055(matchingBytes[3055]),
.io_matchingBytes_3056(matchingBytes[3056]),
.io_matchingBytes_3057(matchingBytes[3057]),
.io_matchingBytes_3058(matchingBytes[3058]),
.io_matchingBytes_3059(matchingBytes[3059]),
.io_matchingBytes_3060(matchingBytes[3060]),
.io_matchingBytes_3061(matchingBytes[3061]),
.io_matchingBytes_3062(matchingBytes[3062]),
.io_matchingBytes_3063(matchingBytes[3063]),
.io_matchingBytes_3064(matchingBytes[3064]),
.io_matchingBytes_3065(matchingBytes[3065]),
.io_matchingBytes_3066(matchingBytes[3066]),
.io_matchingBytes_3067(matchingBytes[3067]),
.io_matchingBytes_3068(matchingBytes[3068]),
.io_matchingBytes_3069(matchingBytes[3069]),
.io_matchingBytes_3070(matchingBytes[3070]),
.io_matchingBytes_3071(matchingBytes[3071]),
.io_matchingBytes_3072(matchingBytes[3072]),
.io_matchingBytes_3073(matchingBytes[3073]),
.io_matchingBytes_3074(matchingBytes[3074]),
.io_matchingBytes_3075(matchingBytes[3075]),
.io_matchingBytes_3076(matchingBytes[3076]),
.io_matchingBytes_3077(matchingBytes[3077]),
.io_matchingBytes_3078(matchingBytes[3078]),
.io_matchingBytes_3079(matchingBytes[3079]),
.io_matchingBytes_3080(matchingBytes[3080]),
.io_matchingBytes_3081(matchingBytes[3081]),
.io_matchingBytes_3082(matchingBytes[3082]),
.io_matchingBytes_3083(matchingBytes[3083]),
.io_matchingBytes_3084(matchingBytes[3084]),
.io_matchingBytes_3085(matchingBytes[3085]),
.io_matchingBytes_3086(matchingBytes[3086]),
.io_matchingBytes_3087(matchingBytes[3087]),
.io_matchingBytes_3088(matchingBytes[3088]),
.io_matchingBytes_3089(matchingBytes[3089]),
.io_matchingBytes_3090(matchingBytes[3090]),
.io_matchingBytes_3091(matchingBytes[3091]),
.io_matchingBytes_3092(matchingBytes[3092]),
.io_matchingBytes_3093(matchingBytes[3093]),
.io_matchingBytes_3094(matchingBytes[3094]),
.io_matchingBytes_3095(matchingBytes[3095]),
.io_matchingBytes_3096(matchingBytes[3096]),
.io_matchingBytes_3097(matchingBytes[3097]),
.io_matchingBytes_3098(matchingBytes[3098]),
.io_matchingBytes_3099(matchingBytes[3099]),
.io_matchingBytes_3100(matchingBytes[3100]),
.io_matchingBytes_3101(matchingBytes[3101]),
.io_matchingBytes_3102(matchingBytes[3102]),
.io_matchingBytes_3103(matchingBytes[3103]),
.io_matchingBytes_3104(matchingBytes[3104]),
.io_matchingBytes_3105(matchingBytes[3105]),
.io_matchingBytes_3106(matchingBytes[3106]),
.io_matchingBytes_3107(matchingBytes[3107]),
.io_matchingBytes_3108(matchingBytes[3108]),
.io_matchingBytes_3109(matchingBytes[3109]),
.io_matchingBytes_3110(matchingBytes[3110]),
.io_matchingBytes_3111(matchingBytes[3111]),
.io_matchingBytes_3112(matchingBytes[3112]),
.io_matchingBytes_3113(matchingBytes[3113]),
.io_matchingBytes_3114(matchingBytes[3114]),
.io_matchingBytes_3115(matchingBytes[3115]),
.io_matchingBytes_3116(matchingBytes[3116]),
.io_matchingBytes_3117(matchingBytes[3117]),
.io_matchingBytes_3118(matchingBytes[3118]),
.io_matchingBytes_3119(matchingBytes[3119]),
.io_matchingBytes_3120(matchingBytes[3120]),
.io_matchingBytes_3121(matchingBytes[3121]),
.io_matchingBytes_3122(matchingBytes[3122]),
.io_matchingBytes_3123(matchingBytes[3123]),
.io_matchingBytes_3124(matchingBytes[3124]),
.io_matchingBytes_3125(matchingBytes[3125]),
.io_matchingBytes_3126(matchingBytes[3126]),
.io_matchingBytes_3127(matchingBytes[3127]),
.io_matchingBytes_3128(matchingBytes[3128]),
.io_matchingBytes_3129(matchingBytes[3129]),
.io_matchingBytes_3130(matchingBytes[3130]),
.io_matchingBytes_3131(matchingBytes[3131]),
.io_matchingBytes_3132(matchingBytes[3132]),
.io_matchingBytes_3133(matchingBytes[3133]),
.io_matchingBytes_3134(matchingBytes[3134]),
.io_matchingBytes_3135(matchingBytes[3135]),
.io_matchingBytes_3136(matchingBytes[3136]),
.io_matchingBytes_3137(matchingBytes[3137]),
.io_matchingBytes_3138(matchingBytes[3138]),
.io_matchingBytes_3139(matchingBytes[3139]),
.io_matchingBytes_3140(matchingBytes[3140]),
.io_matchingBytes_3141(matchingBytes[3141]),
.io_matchingBytes_3142(matchingBytes[3142]),
.io_matchingBytes_3143(matchingBytes[3143]),
.io_matchingBytes_3144(matchingBytes[3144]),
.io_matchingBytes_3145(matchingBytes[3145]),
.io_matchingBytes_3146(matchingBytes[3146]),
.io_matchingBytes_3147(matchingBytes[3147]),
.io_matchingBytes_3148(matchingBytes[3148]),
.io_matchingBytes_3149(matchingBytes[3149]),
.io_matchingBytes_3150(matchingBytes[3150]),
.io_matchingBytes_3151(matchingBytes[3151]),
.io_matchingBytes_3152(matchingBytes[3152]),
.io_matchingBytes_3153(matchingBytes[3153]),
.io_matchingBytes_3154(matchingBytes[3154]),
.io_matchingBytes_3155(matchingBytes[3155]),
.io_matchingBytes_3156(matchingBytes[3156]),
.io_matchingBytes_3157(matchingBytes[3157]),
.io_matchingBytes_3158(matchingBytes[3158]),
.io_matchingBytes_3159(matchingBytes[3159]),
.io_matchingBytes_3160(matchingBytes[3160]),
.io_matchingBytes_3161(matchingBytes[3161]),
.io_matchingBytes_3162(matchingBytes[3162]),
.io_matchingBytes_3163(matchingBytes[3163]),
.io_matchingBytes_3164(matchingBytes[3164]),
.io_matchingBytes_3165(matchingBytes[3165]),
.io_matchingBytes_3166(matchingBytes[3166]),
.io_matchingBytes_3167(matchingBytes[3167]),
.io_matchingBytes_3168(matchingBytes[3168]),
.io_matchingBytes_3169(matchingBytes[3169]),
.io_matchingBytes_3170(matchingBytes[3170]),
.io_matchingBytes_3171(matchingBytes[3171]),
.io_matchingBytes_3172(matchingBytes[3172]),
.io_matchingBytes_3173(matchingBytes[3173]),
.io_matchingBytes_3174(matchingBytes[3174]),
.io_matchingBytes_3175(matchingBytes[3175]),
.io_matchingBytes_3176(matchingBytes[3176]),
.io_matchingBytes_3177(matchingBytes[3177]),
.io_matchingBytes_3178(matchingBytes[3178]),
.io_matchingBytes_3179(matchingBytes[3179]),
.io_matchingBytes_3180(matchingBytes[3180]),
.io_matchingBytes_3181(matchingBytes[3181]),
.io_matchingBytes_3182(matchingBytes[3182]),
.io_matchingBytes_3183(matchingBytes[3183]),
.io_matchingBytes_3184(matchingBytes[3184]),
.io_matchingBytes_3185(matchingBytes[3185]),
.io_matchingBytes_3186(matchingBytes[3186]),
.io_matchingBytes_3187(matchingBytes[3187]),
.io_matchingBytes_3188(matchingBytes[3188]),
.io_matchingBytes_3189(matchingBytes[3189]),
.io_matchingBytes_3190(matchingBytes[3190]),
.io_matchingBytes_3191(matchingBytes[3191]),
.io_matchingBytes_3192(matchingBytes[3192]),
.io_matchingBytes_3193(matchingBytes[3193]),
.io_matchingBytes_3194(matchingBytes[3194]),
.io_matchingBytes_3195(matchingBytes[3195]),
.io_matchingBytes_3196(matchingBytes[3196]),
.io_matchingBytes_3197(matchingBytes[3197]),
.io_matchingBytes_3198(matchingBytes[3198]),
.io_matchingBytes_3199(matchingBytes[3199]),
.io_matchingBytes_3200(matchingBytes[3200]),
.io_matchingBytes_3201(matchingBytes[3201]),
.io_matchingBytes_3202(matchingBytes[3202]),
.io_matchingBytes_3203(matchingBytes[3203]),
.io_matchingBytes_3204(matchingBytes[3204]),
.io_matchingBytes_3205(matchingBytes[3205]),
.io_matchingBytes_3206(matchingBytes[3206]),
.io_matchingBytes_3207(matchingBytes[3207]),
.io_matchingBytes_3208(matchingBytes[3208]),
.io_matchingBytes_3209(matchingBytes[3209]),
.io_matchingBytes_3210(matchingBytes[3210]),
.io_matchingBytes_3211(matchingBytes[3211]),
.io_matchingBytes_3212(matchingBytes[3212]),
.io_matchingBytes_3213(matchingBytes[3213]),
.io_matchingBytes_3214(matchingBytes[3214]),
.io_matchingBytes_3215(matchingBytes[3215]),
.io_matchingBytes_3216(matchingBytes[3216]),
.io_matchingBytes_3217(matchingBytes[3217]),
.io_matchingBytes_3218(matchingBytes[3218]),
.io_matchingBytes_3219(matchingBytes[3219]),
.io_matchingBytes_3220(matchingBytes[3220]),
.io_matchingBytes_3221(matchingBytes[3221]),
.io_matchingBytes_3222(matchingBytes[3222]),
.io_matchingBytes_3223(matchingBytes[3223]),
.io_matchingBytes_3224(matchingBytes[3224]),
.io_matchingBytes_3225(matchingBytes[3225]),
.io_matchingBytes_3226(matchingBytes[3226]),
.io_matchingBytes_3227(matchingBytes[3227]),
.io_matchingBytes_3228(matchingBytes[3228]),
.io_matchingBytes_3229(matchingBytes[3229]),
.io_matchingBytes_3230(matchingBytes[3230]),
.io_matchingBytes_3231(matchingBytes[3231]),
.io_matchingBytes_3232(matchingBytes[3232]),
.io_matchingBytes_3233(matchingBytes[3233]),
.io_matchingBytes_3234(matchingBytes[3234]),
.io_matchingBytes_3235(matchingBytes[3235]),
.io_matchingBytes_3236(matchingBytes[3236]),
.io_matchingBytes_3237(matchingBytes[3237]),
.io_matchingBytes_3238(matchingBytes[3238]),
.io_matchingBytes_3239(matchingBytes[3239]),
.io_matchingBytes_3240(matchingBytes[3240]),
.io_matchingBytes_3241(matchingBytes[3241]),
.io_matchingBytes_3242(matchingBytes[3242]),
.io_matchingBytes_3243(matchingBytes[3243]),
.io_matchingBytes_3244(matchingBytes[3244]),
.io_matchingBytes_3245(matchingBytes[3245]),
.io_matchingBytes_3246(matchingBytes[3246]),
.io_matchingBytes_3247(matchingBytes[3247]),
.io_matchingBytes_3248(matchingBytes[3248]),
.io_matchingBytes_3249(matchingBytes[3249]),
.io_matchingBytes_3250(matchingBytes[3250]),
.io_matchingBytes_3251(matchingBytes[3251]),
.io_matchingBytes_3252(matchingBytes[3252]),
.io_matchingBytes_3253(matchingBytes[3253]),
.io_matchingBytes_3254(matchingBytes[3254]),
.io_matchingBytes_3255(matchingBytes[3255]),
.io_matchingBytes_3256(matchingBytes[3256]),
.io_matchingBytes_3257(matchingBytes[3257]),
.io_matchingBytes_3258(matchingBytes[3258]),
.io_matchingBytes_3259(matchingBytes[3259]),
.io_matchingBytes_3260(matchingBytes[3260]),
.io_matchingBytes_3261(matchingBytes[3261]),
.io_matchingBytes_3262(matchingBytes[3262]),
.io_matchingBytes_3263(matchingBytes[3263]),
.io_matchingBytes_3264(matchingBytes[3264]),
.io_matchingBytes_3265(matchingBytes[3265]),
.io_matchingBytes_3266(matchingBytes[3266]),
.io_matchingBytes_3267(matchingBytes[3267]),
.io_matchingBytes_3268(matchingBytes[3268]),
.io_matchingBytes_3269(matchingBytes[3269]),
.io_matchingBytes_3270(matchingBytes[3270]),
.io_matchingBytes_3271(matchingBytes[3271]),
.io_matchingBytes_3272(matchingBytes[3272]),
.io_matchingBytes_3273(matchingBytes[3273]),
.io_matchingBytes_3274(matchingBytes[3274]),
.io_matchingBytes_3275(matchingBytes[3275]),
.io_matchingBytes_3276(matchingBytes[3276]),
.io_matchingBytes_3277(matchingBytes[3277]),
.io_matchingBytes_3278(matchingBytes[3278]),
.io_matchingBytes_3279(matchingBytes[3279]),
.io_matchingBytes_3280(matchingBytes[3280]),
.io_matchingBytes_3281(matchingBytes[3281]),
.io_matchingBytes_3282(matchingBytes[3282]),
.io_matchingBytes_3283(matchingBytes[3283]),
.io_matchingBytes_3284(matchingBytes[3284]),
.io_matchingBytes_3285(matchingBytes[3285]),
.io_matchingBytes_3286(matchingBytes[3286]),
.io_matchingBytes_3287(matchingBytes[3287]),
.io_matchingBytes_3288(matchingBytes[3288]),
.io_matchingBytes_3289(matchingBytes[3289]),
.io_matchingBytes_3290(matchingBytes[3290]),
.io_matchingBytes_3291(matchingBytes[3291]),
.io_matchingBytes_3292(matchingBytes[3292]),
.io_matchingBytes_3293(matchingBytes[3293]),
.io_matchingBytes_3294(matchingBytes[3294]),
.io_matchingBytes_3295(matchingBytes[3295]),
.io_matchingBytes_3296(matchingBytes[3296]),
.io_matchingBytes_3297(matchingBytes[3297]),
.io_matchingBytes_3298(matchingBytes[3298]),
.io_matchingBytes_3299(matchingBytes[3299]),
.io_matchingBytes_3300(matchingBytes[3300]),
.io_matchingBytes_3301(matchingBytes[3301]),
.io_matchingBytes_3302(matchingBytes[3302]),
.io_matchingBytes_3303(matchingBytes[3303]),
.io_matchingBytes_3304(matchingBytes[3304]),
.io_matchingBytes_3305(matchingBytes[3305]),
.io_matchingBytes_3306(matchingBytes[3306]),
.io_matchingBytes_3307(matchingBytes[3307]),
.io_matchingBytes_3308(matchingBytes[3308]),
.io_matchingBytes_3309(matchingBytes[3309]),
.io_matchingBytes_3310(matchingBytes[3310]),
.io_matchingBytes_3311(matchingBytes[3311]),
.io_matchingBytes_3312(matchingBytes[3312]),
.io_matchingBytes_3313(matchingBytes[3313]),
.io_matchingBytes_3314(matchingBytes[3314]),
.io_matchingBytes_3315(matchingBytes[3315]),
.io_matchingBytes_3316(matchingBytes[3316]),
.io_matchingBytes_3317(matchingBytes[3317]),
.io_matchingBytes_3318(matchingBytes[3318]),
.io_matchingBytes_3319(matchingBytes[3319]),
.io_matchingBytes_3320(matchingBytes[3320]),
.io_matchingBytes_3321(matchingBytes[3321]),
.io_matchingBytes_3322(matchingBytes[3322]),
.io_matchingBytes_3323(matchingBytes[3323]),
.io_matchingBytes_3324(matchingBytes[3324]),
.io_matchingBytes_3325(matchingBytes[3325]),
.io_matchingBytes_3326(matchingBytes[3326]),
.io_matchingBytes_3327(matchingBytes[3327]),
.io_matchingBytes_3328(matchingBytes[3328]),
.io_matchingBytes_3329(matchingBytes[3329]),
.io_matchingBytes_3330(matchingBytes[3330]),
.io_matchingBytes_3331(matchingBytes[3331]),
.io_matchingBytes_3332(matchingBytes[3332]),
.io_matchingBytes_3333(matchingBytes[3333]),
.io_matchingBytes_3334(matchingBytes[3334]),
.io_matchingBytes_3335(matchingBytes[3335]),
.io_matchingBytes_3336(matchingBytes[3336]),
.io_matchingBytes_3337(matchingBytes[3337]),
.io_matchingBytes_3338(matchingBytes[3338]),
.io_matchingBytes_3339(matchingBytes[3339]),
.io_matchingBytes_3340(matchingBytes[3340]),
.io_matchingBytes_3341(matchingBytes[3341]),
.io_matchingBytes_3342(matchingBytes[3342]),
.io_matchingBytes_3343(matchingBytes[3343]),
.io_matchingBytes_3344(matchingBytes[3344]),
.io_matchingBytes_3345(matchingBytes[3345]),
.io_matchingBytes_3346(matchingBytes[3346]),
.io_matchingBytes_3347(matchingBytes[3347]),
.io_matchingBytes_3348(matchingBytes[3348]),
.io_matchingBytes_3349(matchingBytes[3349]),
.io_matchingBytes_3350(matchingBytes[3350]),
.io_matchingBytes_3351(matchingBytes[3351]),
.io_matchingBytes_3352(matchingBytes[3352]),
.io_matchingBytes_3353(matchingBytes[3353]),
.io_matchingBytes_3354(matchingBytes[3354]),
.io_matchingBytes_3355(matchingBytes[3355]),
.io_matchingBytes_3356(matchingBytes[3356]),
.io_matchingBytes_3357(matchingBytes[3357]),
.io_matchingBytes_3358(matchingBytes[3358]),
.io_matchingBytes_3359(matchingBytes[3359]),
.io_matchingBytes_3360(matchingBytes[3360]),
.io_matchingBytes_3361(matchingBytes[3361]),
.io_matchingBytes_3362(matchingBytes[3362]),
.io_matchingBytes_3363(matchingBytes[3363]),
.io_matchingBytes_3364(matchingBytes[3364]),
.io_matchingBytes_3365(matchingBytes[3365]),
.io_matchingBytes_3366(matchingBytes[3366]),
.io_matchingBytes_3367(matchingBytes[3367]),
.io_matchingBytes_3368(matchingBytes[3368]),
.io_matchingBytes_3369(matchingBytes[3369]),
.io_matchingBytes_3370(matchingBytes[3370]),
.io_matchingBytes_3371(matchingBytes[3371]),
.io_matchingBytes_3372(matchingBytes[3372]),
.io_matchingBytes_3373(matchingBytes[3373]),
.io_matchingBytes_3374(matchingBytes[3374]),
.io_matchingBytes_3375(matchingBytes[3375]),
.io_matchingBytes_3376(matchingBytes[3376]),
.io_matchingBytes_3377(matchingBytes[3377]),
.io_matchingBytes_3378(matchingBytes[3378]),
.io_matchingBytes_3379(matchingBytes[3379]),
.io_matchingBytes_3380(matchingBytes[3380]),
.io_matchingBytes_3381(matchingBytes[3381]),
.io_matchingBytes_3382(matchingBytes[3382]),
.io_matchingBytes_3383(matchingBytes[3383]),
.io_matchingBytes_3384(matchingBytes[3384]),
.io_matchingBytes_3385(matchingBytes[3385]),
.io_matchingBytes_3386(matchingBytes[3386]),
.io_matchingBytes_3387(matchingBytes[3387]),
.io_matchingBytes_3388(matchingBytes[3388]),
.io_matchingBytes_3389(matchingBytes[3389]),
.io_matchingBytes_3390(matchingBytes[3390]),
.io_matchingBytes_3391(matchingBytes[3391]),
.io_matchingBytes_3392(matchingBytes[3392]),
.io_matchingBytes_3393(matchingBytes[3393]),
.io_matchingBytes_3394(matchingBytes[3394]),
.io_matchingBytes_3395(matchingBytes[3395]),
.io_matchingBytes_3396(matchingBytes[3396]),
.io_matchingBytes_3397(matchingBytes[3397]),
.io_matchingBytes_3398(matchingBytes[3398]),
.io_matchingBytes_3399(matchingBytes[3399]),
.io_matchingBytes_3400(matchingBytes[3400]),
.io_matchingBytes_3401(matchingBytes[3401]),
.io_matchingBytes_3402(matchingBytes[3402]),
.io_matchingBytes_3403(matchingBytes[3403]),
.io_matchingBytes_3404(matchingBytes[3404]),
.io_matchingBytes_3405(matchingBytes[3405]),
.io_matchingBytes_3406(matchingBytes[3406]),
.io_matchingBytes_3407(matchingBytes[3407]),
.io_matchingBytes_3408(matchingBytes[3408]),
.io_matchingBytes_3409(matchingBytes[3409]),
.io_matchingBytes_3410(matchingBytes[3410]),
.io_matchingBytes_3411(matchingBytes[3411]),
.io_matchingBytes_3412(matchingBytes[3412]),
.io_matchingBytes_3413(matchingBytes[3413]),
.io_matchingBytes_3414(matchingBytes[3414]),
.io_matchingBytes_3415(matchingBytes[3415]),
.io_matchingBytes_3416(matchingBytes[3416]),
.io_matchingBytes_3417(matchingBytes[3417]),
.io_matchingBytes_3418(matchingBytes[3418]),
.io_matchingBytes_3419(matchingBytes[3419]),
.io_matchingBytes_3420(matchingBytes[3420]),
.io_matchingBytes_3421(matchingBytes[3421]),
.io_matchingBytes_3422(matchingBytes[3422]),
.io_matchingBytes_3423(matchingBytes[3423]),
.io_matchingBytes_3424(matchingBytes[3424]),
.io_matchingBytes_3425(matchingBytes[3425]),
.io_matchingBytes_3426(matchingBytes[3426]),
.io_matchingBytes_3427(matchingBytes[3427]),
.io_matchingBytes_3428(matchingBytes[3428]),
.io_matchingBytes_3429(matchingBytes[3429]),
.io_matchingBytes_3430(matchingBytes[3430]),
.io_matchingBytes_3431(matchingBytes[3431]),
.io_matchingBytes_3432(matchingBytes[3432]),
.io_matchingBytes_3433(matchingBytes[3433]),
.io_matchingBytes_3434(matchingBytes[3434]),
.io_matchingBytes_3435(matchingBytes[3435]),
.io_matchingBytes_3436(matchingBytes[3436]),
.io_matchingBytes_3437(matchingBytes[3437]),
.io_matchingBytes_3438(matchingBytes[3438]),
.io_matchingBytes_3439(matchingBytes[3439]),
.io_matchingBytes_3440(matchingBytes[3440]),
.io_matchingBytes_3441(matchingBytes[3441]),
.io_matchingBytes_3442(matchingBytes[3442]),
.io_matchingBytes_3443(matchingBytes[3443]),
.io_matchingBytes_3444(matchingBytes[3444]),
.io_matchingBytes_3445(matchingBytes[3445]),
.io_matchingBytes_3446(matchingBytes[3446]),
.io_matchingBytes_3447(matchingBytes[3447]),
.io_matchingBytes_3448(matchingBytes[3448]),
.io_matchingBytes_3449(matchingBytes[3449]),
.io_matchingBytes_3450(matchingBytes[3450]),
.io_matchingBytes_3451(matchingBytes[3451]),
.io_matchingBytes_3452(matchingBytes[3452]),
.io_matchingBytes_3453(matchingBytes[3453]),
.io_matchingBytes_3454(matchingBytes[3454]),
.io_matchingBytes_3455(matchingBytes[3455]),
.io_matchingBytes_3456(matchingBytes[3456]),
.io_matchingBytes_3457(matchingBytes[3457]),
.io_matchingBytes_3458(matchingBytes[3458]),
.io_matchingBytes_3459(matchingBytes[3459]),
.io_matchingBytes_3460(matchingBytes[3460]),
.io_matchingBytes_3461(matchingBytes[3461]),
.io_matchingBytes_3462(matchingBytes[3462]),
.io_matchingBytes_3463(matchingBytes[3463]),
.io_matchingBytes_3464(matchingBytes[3464]),
.io_matchingBytes_3465(matchingBytes[3465]),
.io_matchingBytes_3466(matchingBytes[3466]),
.io_matchingBytes_3467(matchingBytes[3467]),
.io_matchingBytes_3468(matchingBytes[3468]),
.io_matchingBytes_3469(matchingBytes[3469]),
.io_matchingBytes_3470(matchingBytes[3470]),
.io_matchingBytes_3471(matchingBytes[3471]),
.io_matchingBytes_3472(matchingBytes[3472]),
.io_matchingBytes_3473(matchingBytes[3473]),
.io_matchingBytes_3474(matchingBytes[3474]),
.io_matchingBytes_3475(matchingBytes[3475]),
.io_matchingBytes_3476(matchingBytes[3476]),
.io_matchingBytes_3477(matchingBytes[3477]),
.io_matchingBytes_3478(matchingBytes[3478]),
.io_matchingBytes_3479(matchingBytes[3479]),
.io_matchingBytes_3480(matchingBytes[3480]),
.io_matchingBytes_3481(matchingBytes[3481]),
.io_matchingBytes_3482(matchingBytes[3482]),
.io_matchingBytes_3483(matchingBytes[3483]),
.io_matchingBytes_3484(matchingBytes[3484]),
.io_matchingBytes_3485(matchingBytes[3485]),
.io_matchingBytes_3486(matchingBytes[3486]),
.io_matchingBytes_3487(matchingBytes[3487]),
.io_matchingBytes_3488(matchingBytes[3488]),
.io_matchingBytes_3489(matchingBytes[3489]),
.io_matchingBytes_3490(matchingBytes[3490]),
.io_matchingBytes_3491(matchingBytes[3491]),
.io_matchingBytes_3492(matchingBytes[3492]),
.io_matchingBytes_3493(matchingBytes[3493]),
.io_matchingBytes_3494(matchingBytes[3494]),
.io_matchingBytes_3495(matchingBytes[3495]),
.io_matchingBytes_3496(matchingBytes[3496]),
.io_matchingBytes_3497(matchingBytes[3497]),
.io_matchingBytes_3498(matchingBytes[3498]),
.io_matchingBytes_3499(matchingBytes[3499]),
.io_matchingBytes_3500(matchingBytes[3500]),
.io_matchingBytes_3501(matchingBytes[3501]),
.io_matchingBytes_3502(matchingBytes[3502]),
.io_matchingBytes_3503(matchingBytes[3503]),
.io_matchingBytes_3504(matchingBytes[3504]),
.io_matchingBytes_3505(matchingBytes[3505]),
.io_matchingBytes_3506(matchingBytes[3506]),
.io_matchingBytes_3507(matchingBytes[3507]),
.io_matchingBytes_3508(matchingBytes[3508]),
.io_matchingBytes_3509(matchingBytes[3509]),
.io_matchingBytes_3510(matchingBytes[3510]),
.io_matchingBytes_3511(matchingBytes[3511]),
.io_matchingBytes_3512(matchingBytes[3512]),
.io_matchingBytes_3513(matchingBytes[3513]),
.io_matchingBytes_3514(matchingBytes[3514]),
.io_matchingBytes_3515(matchingBytes[3515]),
.io_matchingBytes_3516(matchingBytes[3516]),
.io_matchingBytes_3517(matchingBytes[3517]),
.io_matchingBytes_3518(matchingBytes[3518]),
.io_matchingBytes_3519(matchingBytes[3519]),
.io_matchingBytes_3520(matchingBytes[3520]),
.io_matchingBytes_3521(matchingBytes[3521]),
.io_matchingBytes_3522(matchingBytes[3522]),
.io_matchingBytes_3523(matchingBytes[3523]),
.io_matchingBytes_3524(matchingBytes[3524]),
.io_matchingBytes_3525(matchingBytes[3525]),
.io_matchingBytes_3526(matchingBytes[3526]),
.io_matchingBytes_3527(matchingBytes[3527]),
.io_matchingBytes_3528(matchingBytes[3528]),
.io_matchingBytes_3529(matchingBytes[3529]),
.io_matchingBytes_3530(matchingBytes[3530]),
.io_matchingBytes_3531(matchingBytes[3531]),
.io_matchingBytes_3532(matchingBytes[3532]),
.io_matchingBytes_3533(matchingBytes[3533]),
.io_matchingBytes_3534(matchingBytes[3534]),
.io_matchingBytes_3535(matchingBytes[3535]),
.io_matchingBytes_3536(matchingBytes[3536]),
.io_matchingBytes_3537(matchingBytes[3537]),
.io_matchingBytes_3538(matchingBytes[3538]),
.io_matchingBytes_3539(matchingBytes[3539]),
.io_matchingBytes_3540(matchingBytes[3540]),
.io_matchingBytes_3541(matchingBytes[3541]),
.io_matchingBytes_3542(matchingBytes[3542]),
.io_matchingBytes_3543(matchingBytes[3543]),
.io_matchingBytes_3544(matchingBytes[3544]),
.io_matchingBytes_3545(matchingBytes[3545]),
.io_matchingBytes_3546(matchingBytes[3546]),
.io_matchingBytes_3547(matchingBytes[3547]),
.io_matchingBytes_3548(matchingBytes[3548]),
.io_matchingBytes_3549(matchingBytes[3549]),
.io_matchingBytes_3550(matchingBytes[3550]),
.io_matchingBytes_3551(matchingBytes[3551]),
.io_matchingBytes_3552(matchingBytes[3552]),
.io_matchingBytes_3553(matchingBytes[3553]),
.io_matchingBytes_3554(matchingBytes[3554]),
.io_matchingBytes_3555(matchingBytes[3555]),
.io_matchingBytes_3556(matchingBytes[3556]),
.io_matchingBytes_3557(matchingBytes[3557]),
.io_matchingBytes_3558(matchingBytes[3558]),
.io_matchingBytes_3559(matchingBytes[3559]),
.io_matchingBytes_3560(matchingBytes[3560]),
.io_matchingBytes_3561(matchingBytes[3561]),
.io_matchingBytes_3562(matchingBytes[3562]),
.io_matchingBytes_3563(matchingBytes[3563]),
.io_matchingBytes_3564(matchingBytes[3564]),
.io_matchingBytes_3565(matchingBytes[3565]),
.io_matchingBytes_3566(matchingBytes[3566]),
.io_matchingBytes_3567(matchingBytes[3567]),
.io_matchingBytes_3568(matchingBytes[3568]),
.io_matchingBytes_3569(matchingBytes[3569]),
.io_matchingBytes_3570(matchingBytes[3570]),
.io_matchingBytes_3571(matchingBytes[3571]),
.io_matchingBytes_3572(matchingBytes[3572]),
.io_matchingBytes_3573(matchingBytes[3573]),
.io_matchingBytes_3574(matchingBytes[3574]),
.io_matchingBytes_3575(matchingBytes[3575]),
.io_matchingBytes_3576(matchingBytes[3576]),
.io_matchingBytes_3577(matchingBytes[3577]),
.io_matchingBytes_3578(matchingBytes[3578]),
.io_matchingBytes_3579(matchingBytes[3579]),
.io_matchingBytes_3580(matchingBytes[3580]),
.io_matchingBytes_3581(matchingBytes[3581]),
.io_matchingBytes_3582(matchingBytes[3582]),
.io_matchingBytes_3583(matchingBytes[3583]),
.io_matchingBytes_3584(matchingBytes[3584]),
.io_matchingBytes_3585(matchingBytes[3585]),
.io_matchingBytes_3586(matchingBytes[3586]),
.io_matchingBytes_3587(matchingBytes[3587]),
.io_matchingBytes_3588(matchingBytes[3588]),
.io_matchingBytes_3589(matchingBytes[3589]),
.io_matchingBytes_3590(matchingBytes[3590]),
.io_matchingBytes_3591(matchingBytes[3591]),
.io_matchingBytes_3592(matchingBytes[3592]),
.io_matchingBytes_3593(matchingBytes[3593]),
.io_matchingBytes_3594(matchingBytes[3594]),
.io_matchingBytes_3595(matchingBytes[3595]),
.io_matchingBytes_3596(matchingBytes[3596]),
.io_matchingBytes_3597(matchingBytes[3597]),
.io_matchingBytes_3598(matchingBytes[3598]),
.io_matchingBytes_3599(matchingBytes[3599]),
.io_matchingBytes_3600(matchingBytes[3600]),
.io_matchingBytes_3601(matchingBytes[3601]),
.io_matchingBytes_3602(matchingBytes[3602]),
.io_matchingBytes_3603(matchingBytes[3603]),
.io_matchingBytes_3604(matchingBytes[3604]),
.io_matchingBytes_3605(matchingBytes[3605]),
.io_matchingBytes_3606(matchingBytes[3606]),
.io_matchingBytes_3607(matchingBytes[3607]),
.io_matchingBytes_3608(matchingBytes[3608]),
.io_matchingBytes_3609(matchingBytes[3609]),
.io_matchingBytes_3610(matchingBytes[3610]),
.io_matchingBytes_3611(matchingBytes[3611]),
.io_matchingBytes_3612(matchingBytes[3612]),
.io_matchingBytes_3613(matchingBytes[3613]),
.io_matchingBytes_3614(matchingBytes[3614]),
.io_matchingBytes_3615(matchingBytes[3615]),
.io_matchingBytes_3616(matchingBytes[3616]),
.io_matchingBytes_3617(matchingBytes[3617]),
.io_matchingBytes_3618(matchingBytes[3618]),
.io_matchingBytes_3619(matchingBytes[3619]),
.io_matchingBytes_3620(matchingBytes[3620]),
.io_matchingBytes_3621(matchingBytes[3621]),
.io_matchingBytes_3622(matchingBytes[3622]),
.io_matchingBytes_3623(matchingBytes[3623]),
.io_matchingBytes_3624(matchingBytes[3624]),
.io_matchingBytes_3625(matchingBytes[3625]),
.io_matchingBytes_3626(matchingBytes[3626]),
.io_matchingBytes_3627(matchingBytes[3627]),
.io_matchingBytes_3628(matchingBytes[3628]),
.io_matchingBytes_3629(matchingBytes[3629]),
.io_matchingBytes_3630(matchingBytes[3630]),
.io_matchingBytes_3631(matchingBytes[3631]),
.io_matchingBytes_3632(matchingBytes[3632]),
.io_matchingBytes_3633(matchingBytes[3633]),
.io_matchingBytes_3634(matchingBytes[3634]),
.io_matchingBytes_3635(matchingBytes[3635]),
.io_matchingBytes_3636(matchingBytes[3636]),
.io_matchingBytes_3637(matchingBytes[3637]),
.io_matchingBytes_3638(matchingBytes[3638]),
.io_matchingBytes_3639(matchingBytes[3639]),
.io_matchingBytes_3640(matchingBytes[3640]),
.io_matchingBytes_3641(matchingBytes[3641]),
.io_matchingBytes_3642(matchingBytes[3642]),
.io_matchingBytes_3643(matchingBytes[3643]),
.io_matchingBytes_3644(matchingBytes[3644]),
.io_matchingBytes_3645(matchingBytes[3645]),
.io_matchingBytes_3646(matchingBytes[3646]),
.io_matchingBytes_3647(matchingBytes[3647]),
.io_matchingBytes_3648(matchingBytes[3648]),
.io_matchingBytes_3649(matchingBytes[3649]),
.io_matchingBytes_3650(matchingBytes[3650]),
.io_matchingBytes_3651(matchingBytes[3651]),
.io_matchingBytes_3652(matchingBytes[3652]),
.io_matchingBytes_3653(matchingBytes[3653]),
.io_matchingBytes_3654(matchingBytes[3654]),
.io_matchingBytes_3655(matchingBytes[3655]),
.io_matchingBytes_3656(matchingBytes[3656]),
.io_matchingBytes_3657(matchingBytes[3657]),
.io_matchingBytes_3658(matchingBytes[3658]),
.io_matchingBytes_3659(matchingBytes[3659]),
.io_matchingBytes_3660(matchingBytes[3660]),
.io_matchingBytes_3661(matchingBytes[3661]),
.io_matchingBytes_3662(matchingBytes[3662]),
.io_matchingBytes_3663(matchingBytes[3663]),
.io_matchingBytes_3664(matchingBytes[3664]),
.io_matchingBytes_3665(matchingBytes[3665]),
.io_matchingBytes_3666(matchingBytes[3666]),
.io_matchingBytes_3667(matchingBytes[3667]),
.io_matchingBytes_3668(matchingBytes[3668]),
.io_matchingBytes_3669(matchingBytes[3669]),
.io_matchingBytes_3670(matchingBytes[3670]),
.io_matchingBytes_3671(matchingBytes[3671]),
.io_matchingBytes_3672(matchingBytes[3672]),
.io_matchingBytes_3673(matchingBytes[3673]),
.io_matchingBytes_3674(matchingBytes[3674]),
.io_matchingBytes_3675(matchingBytes[3675]),
.io_matchingBytes_3676(matchingBytes[3676]),
.io_matchingBytes_3677(matchingBytes[3677]),
.io_matchingBytes_3678(matchingBytes[3678]),
.io_matchingBytes_3679(matchingBytes[3679]),
.io_matchingBytes_3680(matchingBytes[3680]),
.io_matchingBytes_3681(matchingBytes[3681]),
.io_matchingBytes_3682(matchingBytes[3682]),
.io_matchingBytes_3683(matchingBytes[3683]),
.io_matchingBytes_3684(matchingBytes[3684]),
.io_matchingBytes_3685(matchingBytes[3685]),
.io_matchingBytes_3686(matchingBytes[3686]),
.io_matchingBytes_3687(matchingBytes[3687]),
.io_matchingBytes_3688(matchingBytes[3688]),
.io_matchingBytes_3689(matchingBytes[3689]),
.io_matchingBytes_3690(matchingBytes[3690]),
.io_matchingBytes_3691(matchingBytes[3691]),
.io_matchingBytes_3692(matchingBytes[3692]),
.io_matchingBytes_3693(matchingBytes[3693]),
.io_matchingBytes_3694(matchingBytes[3694]),
.io_matchingBytes_3695(matchingBytes[3695]),
.io_matchingBytes_3696(matchingBytes[3696]),
.io_matchingBytes_3697(matchingBytes[3697]),
.io_matchingBytes_3698(matchingBytes[3698]),
.io_matchingBytes_3699(matchingBytes[3699]),
.io_matchingBytes_3700(matchingBytes[3700]),
.io_matchingBytes_3701(matchingBytes[3701]),
.io_matchingBytes_3702(matchingBytes[3702]),
.io_matchingBytes_3703(matchingBytes[3703]),
.io_matchingBytes_3704(matchingBytes[3704]),
.io_matchingBytes_3705(matchingBytes[3705]),
.io_matchingBytes_3706(matchingBytes[3706]),
.io_matchingBytes_3707(matchingBytes[3707]),
.io_matchingBytes_3708(matchingBytes[3708]),
.io_matchingBytes_3709(matchingBytes[3709]),
.io_matchingBytes_3710(matchingBytes[3710]),
.io_matchingBytes_3711(matchingBytes[3711]),
.io_matchingBytes_3712(matchingBytes[3712]),
.io_matchingBytes_3713(matchingBytes[3713]),
.io_matchingBytes_3714(matchingBytes[3714]),
.io_matchingBytes_3715(matchingBytes[3715]),
.io_matchingBytes_3716(matchingBytes[3716]),
.io_matchingBytes_3717(matchingBytes[3717]),
.io_matchingBytes_3718(matchingBytes[3718]),
.io_matchingBytes_3719(matchingBytes[3719]),
.io_matchingBytes_3720(matchingBytes[3720]),
.io_matchingBytes_3721(matchingBytes[3721]),
.io_matchingBytes_3722(matchingBytes[3722]),
.io_matchingBytes_3723(matchingBytes[3723]),
.io_matchingBytes_3724(matchingBytes[3724]),
.io_matchingBytes_3725(matchingBytes[3725]),
.io_matchingBytes_3726(matchingBytes[3726]),
.io_matchingBytes_3727(matchingBytes[3727]),
.io_matchingBytes_3728(matchingBytes[3728]),
.io_matchingBytes_3729(matchingBytes[3729]),
.io_matchingBytes_3730(matchingBytes[3730]),
.io_matchingBytes_3731(matchingBytes[3731]),
.io_matchingBytes_3732(matchingBytes[3732]),
.io_matchingBytes_3733(matchingBytes[3733]),
.io_matchingBytes_3734(matchingBytes[3734]),
.io_matchingBytes_3735(matchingBytes[3735]),
.io_matchingBytes_3736(matchingBytes[3736]),
.io_matchingBytes_3737(matchingBytes[3737]),
.io_matchingBytes_3738(matchingBytes[3738]),
.io_matchingBytes_3739(matchingBytes[3739]),
.io_matchingBytes_3740(matchingBytes[3740]),
.io_matchingBytes_3741(matchingBytes[3741]),
.io_matchingBytes_3742(matchingBytes[3742]),
.io_matchingBytes_3743(matchingBytes[3743]),
.io_matchingBytes_3744(matchingBytes[3744]),
.io_matchingBytes_3745(matchingBytes[3745]),
.io_matchingBytes_3746(matchingBytes[3746]),
.io_matchingBytes_3747(matchingBytes[3747]),
.io_matchingBytes_3748(matchingBytes[3748]),
.io_matchingBytes_3749(matchingBytes[3749]),
.io_matchingBytes_3750(matchingBytes[3750]),
.io_matchingBytes_3751(matchingBytes[3751]),
.io_matchingBytes_3752(matchingBytes[3752]),
.io_matchingBytes_3753(matchingBytes[3753]),
.io_matchingBytes_3754(matchingBytes[3754]),
.io_matchingBytes_3755(matchingBytes[3755]),
.io_matchingBytes_3756(matchingBytes[3756]),
.io_matchingBytes_3757(matchingBytes[3757]),
.io_matchingBytes_3758(matchingBytes[3758]),
.io_matchingBytes_3759(matchingBytes[3759]),
.io_matchingBytes_3760(matchingBytes[3760]),
.io_matchingBytes_3761(matchingBytes[3761]),
.io_matchingBytes_3762(matchingBytes[3762]),
.io_matchingBytes_3763(matchingBytes[3763]),
.io_matchingBytes_3764(matchingBytes[3764]),
.io_matchingBytes_3765(matchingBytes[3765]),
.io_matchingBytes_3766(matchingBytes[3766]),
.io_matchingBytes_3767(matchingBytes[3767]),
.io_matchingBytes_3768(matchingBytes[3768]),
.io_matchingBytes_3769(matchingBytes[3769]),
.io_matchingBytes_3770(matchingBytes[3770]),
.io_matchingBytes_3771(matchingBytes[3771]),
.io_matchingBytes_3772(matchingBytes[3772]),
.io_matchingBytes_3773(matchingBytes[3773]),
.io_matchingBytes_3774(matchingBytes[3774]),
.io_matchingBytes_3775(matchingBytes[3775]),
.io_matchingBytes_3776(matchingBytes[3776]),
.io_matchingBytes_3777(matchingBytes[3777]),
.io_matchingBytes_3778(matchingBytes[3778]),
.io_matchingBytes_3779(matchingBytes[3779]),
.io_matchingBytes_3780(matchingBytes[3780]),
.io_matchingBytes_3781(matchingBytes[3781]),
.io_matchingBytes_3782(matchingBytes[3782]),
.io_matchingBytes_3783(matchingBytes[3783]),
.io_matchingBytes_3784(matchingBytes[3784]),
.io_matchingBytes_3785(matchingBytes[3785]),
.io_matchingBytes_3786(matchingBytes[3786]),
.io_matchingBytes_3787(matchingBytes[3787]),
.io_matchingBytes_3788(matchingBytes[3788]),
.io_matchingBytes_3789(matchingBytes[3789]),
.io_matchingBytes_3790(matchingBytes[3790]),
.io_matchingBytes_3791(matchingBytes[3791]),
.io_matchingBytes_3792(matchingBytes[3792]),
.io_matchingBytes_3793(matchingBytes[3793]),
.io_matchingBytes_3794(matchingBytes[3794]),
.io_matchingBytes_3795(matchingBytes[3795]),
.io_matchingBytes_3796(matchingBytes[3796]),
.io_matchingBytes_3797(matchingBytes[3797]),
.io_matchingBytes_3798(matchingBytes[3798]),
.io_matchingBytes_3799(matchingBytes[3799]),
.io_matchingBytes_3800(matchingBytes[3800]),
.io_matchingBytes_3801(matchingBytes[3801]),
.io_matchingBytes_3802(matchingBytes[3802]),
.io_matchingBytes_3803(matchingBytes[3803]),
.io_matchingBytes_3804(matchingBytes[3804]),
.io_matchingBytes_3805(matchingBytes[3805]),
.io_matchingBytes_3806(matchingBytes[3806]),
.io_matchingBytes_3807(matchingBytes[3807]),
.io_matchingBytes_3808(matchingBytes[3808]),
.io_matchingBytes_3809(matchingBytes[3809]),
.io_matchingBytes_3810(matchingBytes[3810]),
.io_matchingBytes_3811(matchingBytes[3811]),
.io_matchingBytes_3812(matchingBytes[3812]),
.io_matchingBytes_3813(matchingBytes[3813]),
.io_matchingBytes_3814(matchingBytes[3814]),
.io_matchingBytes_3815(matchingBytes[3815]),
.io_matchingBytes_3816(matchingBytes[3816]),
.io_matchingBytes_3817(matchingBytes[3817]),
.io_matchingBytes_3818(matchingBytes[3818]),
.io_matchingBytes_3819(matchingBytes[3819]),
.io_matchingBytes_3820(matchingBytes[3820]),
.io_matchingBytes_3821(matchingBytes[3821]),
.io_matchingBytes_3822(matchingBytes[3822]),
.io_matchingBytes_3823(matchingBytes[3823]),
.io_matchingBytes_3824(matchingBytes[3824]),
.io_matchingBytes_3825(matchingBytes[3825]),
.io_matchingBytes_3826(matchingBytes[3826]),
.io_matchingBytes_3827(matchingBytes[3827]),
.io_matchingBytes_3828(matchingBytes[3828]),
.io_matchingBytes_3829(matchingBytes[3829]),
.io_matchingBytes_3830(matchingBytes[3830]),
.io_matchingBytes_3831(matchingBytes[3831]),
.io_matchingBytes_3832(matchingBytes[3832]),
.io_matchingBytes_3833(matchingBytes[3833]),
.io_matchingBytes_3834(matchingBytes[3834]),
.io_matchingBytes_3835(matchingBytes[3835]),
.io_matchingBytes_3836(matchingBytes[3836]),
.io_matchingBytes_3837(matchingBytes[3837]),
.io_matchingBytes_3838(matchingBytes[3838]),
.io_matchingBytes_3839(matchingBytes[3839]),
.io_matchingBytes_3840(matchingBytes[3840]),
.io_matchingBytes_3841(matchingBytes[3841]),
.io_matchingBytes_3842(matchingBytes[3842]),
.io_matchingBytes_3843(matchingBytes[3843]),
.io_matchingBytes_3844(matchingBytes[3844]),
.io_matchingBytes_3845(matchingBytes[3845]),
.io_matchingBytes_3846(matchingBytes[3846]),
.io_matchingBytes_3847(matchingBytes[3847]),
.io_matchingBytes_3848(matchingBytes[3848]),
.io_matchingBytes_3849(matchingBytes[3849]),
.io_matchingBytes_3850(matchingBytes[3850]),
.io_matchingBytes_3851(matchingBytes[3851]),
.io_matchingBytes_3852(matchingBytes[3852]),
.io_matchingBytes_3853(matchingBytes[3853]),
.io_matchingBytes_3854(matchingBytes[3854]),
.io_matchingBytes_3855(matchingBytes[3855]),
.io_matchingBytes_3856(matchingBytes[3856]),
.io_matchingBytes_3857(matchingBytes[3857]),
.io_matchingBytes_3858(matchingBytes[3858]),
.io_matchingBytes_3859(matchingBytes[3859]),
.io_matchingBytes_3860(matchingBytes[3860]),
.io_matchingBytes_3861(matchingBytes[3861]),
.io_matchingBytes_3862(matchingBytes[3862]),
.io_matchingBytes_3863(matchingBytes[3863]),
.io_matchingBytes_3864(matchingBytes[3864]),
.io_matchingBytes_3865(matchingBytes[3865]),
.io_matchingBytes_3866(matchingBytes[3866]),
.io_matchingBytes_3867(matchingBytes[3867]),
.io_matchingBytes_3868(matchingBytes[3868]),
.io_matchingBytes_3869(matchingBytes[3869]),
.io_matchingBytes_3870(matchingBytes[3870]),
.io_matchingBytes_3871(matchingBytes[3871]),
.io_matchingBytes_3872(matchingBytes[3872]),
.io_matchingBytes_3873(matchingBytes[3873]),
.io_matchingBytes_3874(matchingBytes[3874]),
.io_matchingBytes_3875(matchingBytes[3875]),
.io_matchingBytes_3876(matchingBytes[3876]),
.io_matchingBytes_3877(matchingBytes[3877]),
.io_matchingBytes_3878(matchingBytes[3878]),
.io_matchingBytes_3879(matchingBytes[3879]),
.io_matchingBytes_3880(matchingBytes[3880]),
.io_matchingBytes_3881(matchingBytes[3881]),
.io_matchingBytes_3882(matchingBytes[3882]),
.io_matchingBytes_3883(matchingBytes[3883]),
.io_matchingBytes_3884(matchingBytes[3884]),
.io_matchingBytes_3885(matchingBytes[3885]),
.io_matchingBytes_3886(matchingBytes[3886]),
.io_matchingBytes_3887(matchingBytes[3887]),
.io_matchingBytes_3888(matchingBytes[3888]),
.io_matchingBytes_3889(matchingBytes[3889]),
.io_matchingBytes_3890(matchingBytes[3890]),
.io_matchingBytes_3891(matchingBytes[3891]),
.io_matchingBytes_3892(matchingBytes[3892]),
.io_matchingBytes_3893(matchingBytes[3893]),
.io_matchingBytes_3894(matchingBytes[3894]),
.io_matchingBytes_3895(matchingBytes[3895]),
.io_matchingBytes_3896(matchingBytes[3896]),
.io_matchingBytes_3897(matchingBytes[3897]),
.io_matchingBytes_3898(matchingBytes[3898]),
.io_matchingBytes_3899(matchingBytes[3899]),
.io_matchingBytes_3900(matchingBytes[3900]),
.io_matchingBytes_3901(matchingBytes[3901]),
.io_matchingBytes_3902(matchingBytes[3902]),
.io_matchingBytes_3903(matchingBytes[3903]),
.io_matchingBytes_3904(matchingBytes[3904]),
.io_matchingBytes_3905(matchingBytes[3905]),
.io_matchingBytes_3906(matchingBytes[3906]),
.io_matchingBytes_3907(matchingBytes[3907]),
.io_matchingBytes_3908(matchingBytes[3908]),
.io_matchingBytes_3909(matchingBytes[3909]),
.io_matchingBytes_3910(matchingBytes[3910]),
.io_matchingBytes_3911(matchingBytes[3911]),
.io_matchingBytes_3912(matchingBytes[3912]),
.io_matchingBytes_3913(matchingBytes[3913]),
.io_matchingBytes_3914(matchingBytes[3914]),
.io_matchingBytes_3915(matchingBytes[3915]),
.io_matchingBytes_3916(matchingBytes[3916]),
.io_matchingBytes_3917(matchingBytes[3917]),
.io_matchingBytes_3918(matchingBytes[3918]),
.io_matchingBytes_3919(matchingBytes[3919]),
.io_matchingBytes_3920(matchingBytes[3920]),
.io_matchingBytes_3921(matchingBytes[3921]),
.io_matchingBytes_3922(matchingBytes[3922]),
.io_matchingBytes_3923(matchingBytes[3923]),
.io_matchingBytes_3924(matchingBytes[3924]),
.io_matchingBytes_3925(matchingBytes[3925]),
.io_matchingBytes_3926(matchingBytes[3926]),
.io_matchingBytes_3927(matchingBytes[3927]),
.io_matchingBytes_3928(matchingBytes[3928]),
.io_matchingBytes_3929(matchingBytes[3929]),
.io_matchingBytes_3930(matchingBytes[3930]),
.io_matchingBytes_3931(matchingBytes[3931]),
.io_matchingBytes_3932(matchingBytes[3932]),
.io_matchingBytes_3933(matchingBytes[3933]),
.io_matchingBytes_3934(matchingBytes[3934]),
.io_matchingBytes_3935(matchingBytes[3935]),
.io_matchingBytes_3936(matchingBytes[3936]),
.io_matchingBytes_3937(matchingBytes[3937]),
.io_matchingBytes_3938(matchingBytes[3938]),
.io_matchingBytes_3939(matchingBytes[3939]),
.io_matchingBytes_3940(matchingBytes[3940]),
.io_matchingBytes_3941(matchingBytes[3941]),
.io_matchingBytes_3942(matchingBytes[3942]),
.io_matchingBytes_3943(matchingBytes[3943]),
.io_matchingBytes_3944(matchingBytes[3944]),
.io_matchingBytes_3945(matchingBytes[3945]),
.io_matchingBytes_3946(matchingBytes[3946]),
.io_matchingBytes_3947(matchingBytes[3947]),
.io_matchingBytes_3948(matchingBytes[3948]),
.io_matchingBytes_3949(matchingBytes[3949]),
.io_matchingBytes_3950(matchingBytes[3950]),
.io_matchingBytes_3951(matchingBytes[3951]),
.io_matchingBytes_3952(matchingBytes[3952]),
.io_matchingBytes_3953(matchingBytes[3953]),
.io_matchingBytes_3954(matchingBytes[3954]),
.io_matchingBytes_3955(matchingBytes[3955]),
.io_matchingBytes_3956(matchingBytes[3956]),
.io_matchingBytes_3957(matchingBytes[3957]),
.io_matchingBytes_3958(matchingBytes[3958]),
.io_matchingBytes_3959(matchingBytes[3959]),
.io_matchingBytes_3960(matchingBytes[3960]),
.io_matchingBytes_3961(matchingBytes[3961]),
.io_matchingBytes_3962(matchingBytes[3962]),
.io_matchingBytes_3963(matchingBytes[3963]),
.io_matchingBytes_3964(matchingBytes[3964]),
.io_matchingBytes_3965(matchingBytes[3965]),
.io_matchingBytes_3966(matchingBytes[3966]),
.io_matchingBytes_3967(matchingBytes[3967]),
.io_matchingBytes_3968(matchingBytes[3968]),
.io_matchingBytes_3969(matchingBytes[3969]),
.io_matchingBytes_3970(matchingBytes[3970]),
.io_matchingBytes_3971(matchingBytes[3971]),
.io_matchingBytes_3972(matchingBytes[3972]),
.io_matchingBytes_3973(matchingBytes[3973]),
.io_matchingBytes_3974(matchingBytes[3974]),
.io_matchingBytes_3975(matchingBytes[3975]),
.io_matchingBytes_3976(matchingBytes[3976]),
.io_matchingBytes_3977(matchingBytes[3977]),
.io_matchingBytes_3978(matchingBytes[3978]),
.io_matchingBytes_3979(matchingBytes[3979]),
.io_matchingBytes_3980(matchingBytes[3980]),
.io_matchingBytes_3981(matchingBytes[3981]),
.io_matchingBytes_3982(matchingBytes[3982]),
.io_matchingBytes_3983(matchingBytes[3983]),
.io_matchingBytes_3984(matchingBytes[3984]),
.io_matchingBytes_3985(matchingBytes[3985]),
.io_matchingBytes_3986(matchingBytes[3986]),
.io_matchingBytes_3987(matchingBytes[3987]),
.io_matchingBytes_3988(matchingBytes[3988]),
.io_matchingBytes_3989(matchingBytes[3989]),
.io_matchingBytes_3990(matchingBytes[3990]),
.io_matchingBytes_3991(matchingBytes[3991]),
.io_matchingBytes_3992(matchingBytes[3992]),
.io_matchingBytes_3993(matchingBytes[3993]),
.io_matchingBytes_3994(matchingBytes[3994]),
.io_matchingBytes_3995(matchingBytes[3995]),
.io_matchingBytes_3996(matchingBytes[3996]),
.io_matchingBytes_3997(matchingBytes[3997]),
.io_matchingBytes_3998(matchingBytes[3998]),
.io_matchingBytes_3999(matchingBytes[3999]),
.io_matchingBytes_4000(matchingBytes[4000]),
.io_matchingBytes_4001(matchingBytes[4001]),
.io_matchingBytes_4002(matchingBytes[4002]),
.io_matchingBytes_4003(matchingBytes[4003]),
.io_matchingBytes_4004(matchingBytes[4004]),
.io_matchingBytes_4005(matchingBytes[4005]),
.io_matchingBytes_4006(matchingBytes[4006]),
.io_matchingBytes_4007(matchingBytes[4007]),
.io_matchingBytes_4008(matchingBytes[4008]),
.io_matchingBytes_4009(matchingBytes[4009]),
.io_matchingBytes_4010(matchingBytes[4010]),
.io_matchingBytes_4011(matchingBytes[4011]),
.io_matchingBytes_4012(matchingBytes[4012]),
.io_matchingBytes_4013(matchingBytes[4013]),
.io_matchingBytes_4014(matchingBytes[4014]),
.io_matchingBytes_4015(matchingBytes[4015]),
.io_matchingBytes_4016(matchingBytes[4016]),
.io_matchingBytes_4017(matchingBytes[4017]),
.io_matchingBytes_4018(matchingBytes[4018]),
.io_matchingBytes_4019(matchingBytes[4019]),
.io_matchingBytes_4020(matchingBytes[4020]),
.io_matchingBytes_4021(matchingBytes[4021]),
.io_matchingBytes_4022(matchingBytes[4022]),
.io_matchingBytes_4023(matchingBytes[4023]),
.io_matchingBytes_4024(matchingBytes[4024]),
.io_matchingBytes_4025(matchingBytes[4025]),
.io_matchingBytes_4026(matchingBytes[4026]),
.io_matchingBytes_4027(matchingBytes[4027]),
.io_matchingBytes_4028(matchingBytes[4028]),
.io_matchingBytes_4029(matchingBytes[4029]),
.io_matchingBytes_4030(matchingBytes[4030]),
.io_matchingBytes_4031(matchingBytes[4031]),
.io_matchingBytes_4032(matchingBytes[4032]),
.io_matchingBytes_4033(matchingBytes[4033]),
.io_matchingBytes_4034(matchingBytes[4034]),
.io_matchingBytes_4035(matchingBytes[4035]),
.io_matchingBytes_4036(matchingBytes[4036]),
.io_matchingBytes_4037(matchingBytes[4037]),
.io_matchingBytes_4038(matchingBytes[4038]),
.io_matchingBytes_4039(matchingBytes[4039]),
.io_matchingBytes_4040(matchingBytes[4040]),
.io_matchingBytes_4041(matchingBytes[4041]),
.io_matchingBytes_4042(matchingBytes[4042]),
.io_matchingBytes_4043(matchingBytes[4043]),
.io_matchingBytes_4044(matchingBytes[4044]),
.io_matchingBytes_4045(matchingBytes[4045]),
.io_matchingBytes_4046(matchingBytes[4046]),
.io_matchingBytes_4047(matchingBytes[4047]),
.io_matchingBytes_4048(matchingBytes[4048]),
.io_matchingBytes_4049(matchingBytes[4049]),
.io_matchingBytes_4050(matchingBytes[4050]),
.io_matchingBytes_4051(matchingBytes[4051]),
.io_matchingBytes_4052(matchingBytes[4052]),
.io_matchingBytes_4053(matchingBytes[4053]),
.io_matchingBytes_4054(matchingBytes[4054]),
.io_matchingBytes_4055(matchingBytes[4055]),
.io_matchingBytes_4056(matchingBytes[4056]),
.io_matchingBytes_4057(matchingBytes[4057]),
.io_matchingBytes_4058(matchingBytes[4058]),
.io_matchingBytes_4059(matchingBytes[4059]),
.io_matchingBytes_4060(matchingBytes[4060]),
.io_matchingBytes_4061(matchingBytes[4061]),
.io_matchingBytes_4062(matchingBytes[4062]),
.io_matchingBytes_4063(matchingBytes[4063]),
.io_matchingBytes_4064(matchingBytes[4064]),
.io_matchingBytes_4065(matchingBytes[4065]),
.io_matchingBytes_4066(matchingBytes[4066]),
.io_matchingBytes_4067(matchingBytes[4067]),
.io_matchingBytes_4068(matchingBytes[4068]),
.io_matchingBytes_4069(matchingBytes[4069]),
.io_matchingBytes_4070(matchingBytes[4070]),
.io_matchingBytes_4071(matchingBytes[4071]),
.io_matchingBytes_4072(matchingBytes[4072]),
.io_matchingBytes_4073(matchingBytes[4073]),
.io_matchingBytes_4074(matchingBytes[4074]),
.io_matchingBytes_4075(matchingBytes[4075]),
.io_matchingBytes_4076(matchingBytes[4076]),
.io_matchingBytes_4077(matchingBytes[4077]),
.io_matchingBytes_4078(matchingBytes[4078]),
.io_matchingBytes_4079(matchingBytes[4079]),
.io_matchingBytes_4080(matchingBytes[4080]),
.io_matchingBytes_4081(matchingBytes[4081]),
.io_matchingBytes_4082(matchingBytes[4082]),
.io_matchingBytes_4083(matchingBytes[4083]),
.io_matchingBytes_4084(matchingBytes[4084]),
.io_matchingBytes_4085(matchingBytes[4085]),
.io_matchingBytes_4086(matchingBytes[4086]),
.io_matchingBytes_4087(matchingBytes[4087]),
.io_matchingBytes_4088(matchingBytes[4088]),
.io_matchingBytes_4089(matchingBytes[4089]),
.io_matchingBytes_4090(matchingBytes[4090]),
.io_matchingBytes_4091(matchingBytes[4091]),
.io_matchingBytes_4092(matchingBytes[4092]),
.io_matchingBytes_4093(matchingBytes[4093]),
.io_matchingBytes_4094(matchingBytes[4094]),
.io_matchingBytes_4095(matchingBytes[4095]),
.io_numberOfMatchingBytes(numberOfMatchingBytes),
.io_lz77CompressedBytes(lz77CompressedBytes),
.io_huffmanCompressedBytes(huffmanCompressedBytes)
);

endmodule

