`timescale 1ns/1ps
module lzwAndHuffmanTestbench();
reg clock, reset, start;
reg [7:0] decompressedDataIn [0:4095];
wire [7:0] decompressedDataOut [0:4095];
wire decompressorFinished;
reg decompressorFinishedPrevious;
integer r, file, fileIterator;
// This is used to determine what data from the testbench input file to read
integer loopCount;
integer desiredLoop = 4;
always @(posedge clock) decompressorFinishedPrevious <= decompressorFinished;

integer count;
integer clockCount;

lzwAndHuffmanWrapper hcdw(
  .clock(clock),
  .reset(reset),
  .start(start),
  .dataIn(decompressedDataIn),
  .dataOut(decompressedDataOut),
  .finished(decompressorFinished)
);

wire inputEqualsOutput;

reg [0:4095] matchByte;
always @(*) begin
  for(count = 0; count < 4096; count = count + 1) begin
    matchByte[count] = decompressedDataIn[count] == decompressedDataOut[count];
  end
end

assign inputEqualsOutput = &matchByte;

initial begin
	$dumpfile("traceOutput.fst");
	$dumpvars(0,lzwAndHuffmanTestbench);
end

initial
  begin
    clock = 0;
    reset = 0;
    start = 0;
    #10;
    $display("testing");
    reset = 1;
    clock = 1;
    #10;
    $display("testing");
    clock = 0;
    #10;
    $display("testing");
    clock = 1;
    #10;
    $display("testing");
    clock = 0;
    #10;
    $display("testing");
    reset = 0;
    $display("testing");
/*
    decompressedDataIn[0] = 127;
    $display("testing");
decompressedDataIn[1] = 69;
    $display("testing");
decompressedDataIn[2] = 76;
    $display("testing");
decompressedDataIn[3] = 70;
    $display("testing");
decompressedDataIn[4] = 2;
    $display("testing");
decompressedDataIn[5] = 1;
    $display("testing");
decompressedDataIn[6] = 1;
    $display("testing");
decompressedDataIn[7] = 0;
    $display("testing");
decompressedDataIn[8] = 0;
    $display("testing");
decompressedDataIn[9] = 0;
    $display("testing");
decompressedDataIn[10] = 0;
    $display("testing");
decompressedDataIn[11] = 0;
    $display("testing");
decompressedDataIn[12] = 0;
    $display("testing");
decompressedDataIn[13] = 0;
decompressedDataIn[14] = 0;
decompressedDataIn[15] = 0;
decompressedDataIn[16] = 4;
decompressedDataIn[17] = 0;
decompressedDataIn[18] = 62;
decompressedDataIn[19] = 0;
decompressedDataIn[20] = 1;
decompressedDataIn[21] = 0;
decompressedDataIn[22] = 0;
decompressedDataIn[23] = 0;
decompressedDataIn[24] = 0;
decompressedDataIn[25] = 0;
decompressedDataIn[26] = 0;
decompressedDataIn[27] = 0;
decompressedDataIn[28] = 0;
decompressedDataIn[29] = 0;
decompressedDataIn[30] = 0;
decompressedDataIn[31] = 0;
decompressedDataIn[32] = 64;
decompressedDataIn[33] = 0;
decompressedDataIn[34] = 0;
decompressedDataIn[35] = 0;
decompressedDataIn[36] = 0;
decompressedDataIn[37] = 0;
decompressedDataIn[38] = 0;
decompressedDataIn[39] = 0;
decompressedDataIn[40] = 32;
decompressedDataIn[41] = 162;
decompressedDataIn[42] = 221;
decompressedDataIn[43] = 23;
decompressedDataIn[44] = 0;
decompressedDataIn[45] = 0;
decompressedDataIn[46] = 0;
decompressedDataIn[47] = 0;
decompressedDataIn[48] = 0;
decompressedDataIn[49] = 0;
decompressedDataIn[50] = 0;
decompressedDataIn[51] = 0;
decompressedDataIn[52] = 64;
decompressedDataIn[53] = 0;
decompressedDataIn[54] = 56;
decompressedDataIn[55] = 0;
decompressedDataIn[56] = 20;
decompressedDataIn[57] = 0;
decompressedDataIn[58] = 64;
decompressedDataIn[59] = 0;
decompressedDataIn[60] = 22;
decompressedDataIn[61] = 0;
decompressedDataIn[62] = 21;
decompressedDataIn[63] = 0;
decompressedDataIn[64] = 4;
decompressedDataIn[65] = 0;
decompressedDataIn[66] = 0;
decompressedDataIn[67] = 0;
decompressedDataIn[68] = 4;
decompressedDataIn[69] = 0;
decompressedDataIn[70] = 0;
decompressedDataIn[71] = 0;
decompressedDataIn[72] = 160;
decompressedDataIn[73] = 4;
decompressedDataIn[74] = 0;
decompressedDataIn[75] = 0;
    $display("testing");
decompressedDataIn[76] = 0;
decompressedDataIn[77] = 0;
decompressedDataIn[78] = 0;
decompressedDataIn[79] = 0;
decompressedDataIn[80] = 0;
decompressedDataIn[81] = 0;
decompressedDataIn[82] = 0;
decompressedDataIn[83] = 0;
decompressedDataIn[84] = 0;
decompressedDataIn[85] = 0;
decompressedDataIn[86] = 0;
decompressedDataIn[87] = 0;
decompressedDataIn[88] = 0;
decompressedDataIn[89] = 0;
decompressedDataIn[90] = 0;
decompressedDataIn[91] = 0;
decompressedDataIn[92] = 0;
decompressedDataIn[93] = 0;
decompressedDataIn[94] = 0;
decompressedDataIn[95] = 0;
decompressedDataIn[96] = 100;
decompressedDataIn[97] = 13;
decompressedDataIn[98] = 0;
decompressedDataIn[99] = 0;
decompressedDataIn[100] = 0;
decompressedDataIn[101] = 0;
decompressedDataIn[102] = 0;
decompressedDataIn[103] = 0;
decompressedDataIn[104] = 0;
decompressedDataIn[105] = 0;
decompressedDataIn[106] = 0;
decompressedDataIn[107] = 0;
decompressedDataIn[108] = 0;
decompressedDataIn[109] = 0;
decompressedDataIn[110] = 0;
decompressedDataIn[111] = 0;
decompressedDataIn[112] = 1;
decompressedDataIn[113] = 0;
decompressedDataIn[114] = 0;
decompressedDataIn[115] = 0;
decompressedDataIn[116] = 0;
decompressedDataIn[117] = 0;
decompressedDataIn[118] = 0;
decompressedDataIn[119] = 0;
decompressedDataIn[120] = 1;
decompressedDataIn[121] = 0;
decompressedDataIn[122] = 0;
decompressedDataIn[123] = 0;
decompressedDataIn[124] = 4;
decompressedDataIn[125] = 0;
decompressedDataIn[126] = 0;
decompressedDataIn[127] = 0;
decompressedDataIn[128] = 4;
decompressedDataIn[129] = 18;
decompressedDataIn[130] = 0;
decompressedDataIn[131] = 0;
decompressedDataIn[132] = 0;
decompressedDataIn[133] = 0;
decompressedDataIn[134] = 0;
decompressedDataIn[135] = 0;
decompressedDataIn[136] = 0;
decompressedDataIn[137] = 32;
decompressedDataIn[138] = 203;
decompressedDataIn[139] = 213;
decompressedDataIn[140] = 109;
decompressedDataIn[141] = 85;
decompressedDataIn[142] = 0;
decompressedDataIn[143] = 0;
decompressedDataIn[144] = 0;
decompressedDataIn[145] = 0;
decompressedDataIn[146] = 0;
decompressedDataIn[147] = 0;
decompressedDataIn[148] = 0;
decompressedDataIn[149] = 0;
decompressedDataIn[150] = 0;
decompressedDataIn[151] = 0;
decompressedDataIn[152] = 0;
decompressedDataIn[153] = 16;
decompressedDataIn[154] = 0;
decompressedDataIn[155] = 0;
decompressedDataIn[156] = 0;
decompressedDataIn[157] = 0;
decompressedDataIn[158] = 0;
decompressedDataIn[159] = 0;
decompressedDataIn[160] = 0;
decompressedDataIn[161] = 16;
decompressedDataIn[162] = 0;
decompressedDataIn[163] = 0;
decompressedDataIn[164] = 0;
decompressedDataIn[165] = 0;
decompressedDataIn[166] = 0;
decompressedDataIn[167] = 0;
decompressedDataIn[168] = 1;
decompressedDataIn[169] = 0;
decompressedDataIn[170] = 0;
decompressedDataIn[171] = 0;
decompressedDataIn[172] = 0;
decompressedDataIn[173] = 0;
decompressedDataIn[174] = 0;
decompressedDataIn[175] = 0;
decompressedDataIn[176] = 1;
decompressedDataIn[177] = 0;
decompressedDataIn[178] = 0;
decompressedDataIn[179] = 0;
decompressedDataIn[180] = 6;
decompressedDataIn[181] = 0;
decompressedDataIn[182] = 0;
decompressedDataIn[183] = 0;
decompressedDataIn[184] = 4;
decompressedDataIn[185] = 34;
decompressedDataIn[186] = 0;
decompressedDataIn[187] = 0;
decompressedDataIn[188] = 0;
decompressedDataIn[189] = 0;
decompressedDataIn[190] = 0;
decompressedDataIn[191] = 0;
decompressedDataIn[192] = 0;
decompressedDataIn[193] = 48;
decompressedDataIn[194] = 203;
decompressedDataIn[195] = 213;
decompressedDataIn[196] = 109;
decompressedDataIn[197] = 85;
decompressedDataIn[198] = 0;
decompressedDataIn[199] = 0;
decompressedDataIn[200] = 0;
decompressedDataIn[201] = 0;
decompressedDataIn[202] = 0;
decompressedDataIn[203] = 0;
decompressedDataIn[204] = 0;
decompressedDataIn[205] = 0;
decompressedDataIn[206] = 0;
decompressedDataIn[207] = 0;
decompressedDataIn[208] = 0;
decompressedDataIn[209] = 16;
decompressedDataIn[210] = 0;
decompressedDataIn[211] = 0;
decompressedDataIn[212] = 0;
decompressedDataIn[213] = 0;
decompressedDataIn[214] = 0;
decompressedDataIn[215] = 0;
decompressedDataIn[216] = 0;
decompressedDataIn[217] = 16;
decompressedDataIn[218] = 0;
decompressedDataIn[219] = 0;
decompressedDataIn[220] = 0;
decompressedDataIn[221] = 0;
decompressedDataIn[222] = 0;
decompressedDataIn[223] = 0;
decompressedDataIn[224] = 1;
decompressedDataIn[225] = 0;
decompressedDataIn[226] = 0;
decompressedDataIn[227] = 0;
decompressedDataIn[228] = 0;
decompressedDataIn[229] = 0;
decompressedDataIn[230] = 0;
decompressedDataIn[231] = 0;
decompressedDataIn[232] = 1;
decompressedDataIn[233] = 0;
decompressedDataIn[234] = 0;
decompressedDataIn[235] = 0;
decompressedDataIn[236] = 6;
decompressedDataIn[237] = 0;
decompressedDataIn[238] = 0;
decompressedDataIn[239] = 0;
decompressedDataIn[240] = 4;
decompressedDataIn[241] = 50;
decompressedDataIn[242] = 0;
decompressedDataIn[243] = 0;
decompressedDataIn[244] = 0;
decompressedDataIn[245] = 0;
decompressedDataIn[246] = 0;
decompressedDataIn[247] = 0;
decompressedDataIn[248] = 0;
decompressedDataIn[249] = 224;
decompressedDataIn[250] = 130;
decompressedDataIn[251] = 215;
decompressedDataIn[252] = 109;
decompressedDataIn[253] = 85;
decompressedDataIn[254] = 0;
decompressedDataIn[255] = 0;
decompressedDataIn[256] = 0;
decompressedDataIn[257] = 0;
decompressedDataIn[258] = 0;
decompressedDataIn[259] = 0;
decompressedDataIn[260] = 0;
decompressedDataIn[261] = 0;
decompressedDataIn[262] = 0;
decompressedDataIn[263] = 0;
decompressedDataIn[264] = 0;
decompressedDataIn[265] = 16;
decompressedDataIn[266] = 2;
decompressedDataIn[267] = 0;
decompressedDataIn[268] = 0;
decompressedDataIn[269] = 0;
decompressedDataIn[270] = 0;
decompressedDataIn[271] = 0;
decompressedDataIn[272] = 0;
decompressedDataIn[273] = 16;
decompressedDataIn[274] = 2;
decompressedDataIn[275] = 0;
    $display("testing");
decompressedDataIn[276] = 0;
decompressedDataIn[277] = 0;
decompressedDataIn[278] = 0;
decompressedDataIn[279] = 0;
decompressedDataIn[280] = 1;
decompressedDataIn[281] = 0;
decompressedDataIn[282] = 0;
decompressedDataIn[283] = 0;
decompressedDataIn[284] = 0;
decompressedDataIn[285] = 0;
decompressedDataIn[286] = 0;
decompressedDataIn[287] = 0;
decompressedDataIn[288] = 1;
decompressedDataIn[289] = 0;
decompressedDataIn[290] = 0;
decompressedDataIn[291] = 0;
decompressedDataIn[292] = 6;
decompressedDataIn[293] = 0;
decompressedDataIn[294] = 0;
decompressedDataIn[295] = 0;
decompressedDataIn[296] = 4;
decompressedDataIn[297] = 66;
decompressedDataIn[298] = 2;
decompressedDataIn[299] = 0;
decompressedDataIn[300] = 0;
decompressedDataIn[301] = 0;
decompressedDataIn[302] = 0;
decompressedDataIn[303] = 0;
decompressedDataIn[304] = 0;
decompressedDataIn[305] = 176;
decompressedDataIn[306] = 31;
decompressedDataIn[307] = 223;
decompressedDataIn[308] = 217;
decompressedDataIn[309] = 127;
decompressedDataIn[310] = 0;
decompressedDataIn[311] = 0;
decompressedDataIn[312] = 0;
decompressedDataIn[313] = 0;
decompressedDataIn[314] = 0;
decompressedDataIn[315] = 0;
decompressedDataIn[316] = 0;
decompressedDataIn[317] = 0;
decompressedDataIn[318] = 0;
decompressedDataIn[319] = 0;
decompressedDataIn[320] = 0;
decompressedDataIn[321] = 144;
decompressedDataIn[322] = 215;
decompressedDataIn[323] = 23;
decompressedDataIn[324] = 0;
decompressedDataIn[325] = 0;
decompressedDataIn[326] = 0;
decompressedDataIn[327] = 0;
decompressedDataIn[328] = 0;
decompressedDataIn[329] = 144;
decompressedDataIn[330] = 215;
decompressedDataIn[331] = 23;
decompressedDataIn[332] = 0;
decompressedDataIn[333] = 0;
decompressedDataIn[334] = 0;
decompressedDataIn[335] = 0;
decompressedDataIn[336] = 1;
decompressedDataIn[337] = 0;
decompressedDataIn[338] = 0;
decompressedDataIn[339] = 0;
decompressedDataIn[340] = 0;
decompressedDataIn[341] = 0;
decompressedDataIn[342] = 0;
decompressedDataIn[343] = 0;
decompressedDataIn[344] = 1;
decompressedDataIn[345] = 0;
decompressedDataIn[346] = 0;
decompressedDataIn[347] = 0;
decompressedDataIn[348] = 4;
decompressedDataIn[349] = 0;
decompressedDataIn[350] = 0;
decompressedDataIn[351] = 0;
decompressedDataIn[352] = 4;
decompressedDataIn[353] = 210;
decompressedDataIn[354] = 217;
decompressedDataIn[355] = 23;
decompressedDataIn[356] = 0;
decompressedDataIn[357] = 0;
decompressedDataIn[358] = 0;
decompressedDataIn[359] = 0;
decompressedDataIn[360] = 0;
decompressedDataIn[361] = 176;
decompressedDataIn[362] = 53;
decompressedDataIn[363] = 247;
decompressedDataIn[364] = 217;
decompressedDataIn[365] = 127;
decompressedDataIn[366] = 0;
decompressedDataIn[367] = 0;
decompressedDataIn[368] = 0;
decompressedDataIn[369] = 0;
decompressedDataIn[370] = 0;
decompressedDataIn[371] = 0;
decompressedDataIn[372] = 0;
decompressedDataIn[373] = 0;
decompressedDataIn[374] = 0;
decompressedDataIn[375] = 0;
decompressedDataIn[376] = 0;
decompressedDataIn[377] = 64;
decompressedDataIn[378] = 0;
decompressedDataIn[379] = 0;
decompressedDataIn[380] = 0;
decompressedDataIn[381] = 0;
decompressedDataIn[382] = 0;
decompressedDataIn[383] = 0;
decompressedDataIn[384] = 0;
decompressedDataIn[385] = 64;
decompressedDataIn[386] = 0;
decompressedDataIn[387] = 0;
decompressedDataIn[388] = 0;
decompressedDataIn[389] = 0;
decompressedDataIn[390] = 0;
decompressedDataIn[391] = 0;
decompressedDataIn[392] = 1;
decompressedDataIn[393] = 0;
decompressedDataIn[394] = 0;
decompressedDataIn[395] = 0;
decompressedDataIn[396] = 0;
decompressedDataIn[397] = 0;
decompressedDataIn[398] = 0;
decompressedDataIn[399] = 0;
decompressedDataIn[400] = 1;
decompressedDataIn[401] = 0;
decompressedDataIn[402] = 0;
decompressedDataIn[403] = 0;
decompressedDataIn[404] = 6;
decompressedDataIn[405] = 0;
decompressedDataIn[406] = 0;
decompressedDataIn[407] = 0;
decompressedDataIn[408] = 4;
decompressedDataIn[409] = 18;
decompressedDataIn[410] = 218;
decompressedDataIn[411] = 23;
decompressedDataIn[412] = 0;
decompressedDataIn[413] = 0;
decompressedDataIn[414] = 0;
decompressedDataIn[415] = 0;
decompressedDataIn[416] = 0;
decompressedDataIn[417] = 240;
decompressedDataIn[418] = 53;
decompressedDataIn[419] = 247;
decompressedDataIn[420] = 217;
decompressedDataIn[421] = 127;
decompressedDataIn[422] = 0;
decompressedDataIn[423] = 0;
decompressedDataIn[424] = 0;
decompressedDataIn[425] = 0;
decompressedDataIn[426] = 0;
decompressedDataIn[427] = 0;
decompressedDataIn[428] = 0;
decompressedDataIn[429] = 0;
decompressedDataIn[430] = 0;
decompressedDataIn[431] = 0;
decompressedDataIn[432] = 0;
decompressedDataIn[433] = 32;
decompressedDataIn[434] = 0;
decompressedDataIn[435] = 0;
decompressedDataIn[436] = 0;
decompressedDataIn[437] = 0;
decompressedDataIn[438] = 0;
decompressedDataIn[439] = 0;
decompressedDataIn[440] = 0;
decompressedDataIn[441] = 32;
decompressedDataIn[442] = 0;
decompressedDataIn[443] = 0;
decompressedDataIn[444] = 0;
decompressedDataIn[445] = 0;
decompressedDataIn[446] = 0;
decompressedDataIn[447] = 0;
decompressedDataIn[448] = 1;
decompressedDataIn[449] = 0;
decompressedDataIn[450] = 0;
decompressedDataIn[451] = 0;
decompressedDataIn[452] = 0;
decompressedDataIn[453] = 0;
decompressedDataIn[454] = 0;
decompressedDataIn[455] = 0;
decompressedDataIn[456] = 1;
decompressedDataIn[457] = 0;
decompressedDataIn[458] = 0;
decompressedDataIn[459] = 0;
decompressedDataIn[460] = 6;
decompressedDataIn[461] = 0;
decompressedDataIn[462] = 0;
decompressedDataIn[463] = 0;
decompressedDataIn[464] = 4;
decompressedDataIn[465] = 50;
decompressedDataIn[466] = 218;
decompressedDataIn[467] = 23;
decompressedDataIn[468] = 0;
decompressedDataIn[469] = 0;
decompressedDataIn[470] = 0;
decompressedDataIn[471] = 0;
decompressedDataIn[472] = 0;
decompressedDataIn[473] = 16;
decompressedDataIn[474] = 54;
decompressedDataIn[475] = 247;
decompressedDataIn[476] = 217;
decompressedDataIn[477] = 127;
decompressedDataIn[478] = 0;
decompressedDataIn[479] = 0;
decompressedDataIn[480] = 0;
decompressedDataIn[481] = 0;
decompressedDataIn[482] = 0;
decompressedDataIn[483] = 0;
decompressedDataIn[484] = 0;
decompressedDataIn[485] = 0;
decompressedDataIn[486] = 0;
decompressedDataIn[487] = 0;
decompressedDataIn[488] = 0;
decompressedDataIn[489] = 64;
decompressedDataIn[490] = 0;
decompressedDataIn[491] = 0;
decompressedDataIn[492] = 0;
decompressedDataIn[493] = 0;
decompressedDataIn[494] = 0;
decompressedDataIn[495] = 0;
decompressedDataIn[496] = 0;
decompressedDataIn[497] = 64;
decompressedDataIn[498] = 0;
decompressedDataIn[499] = 0;
decompressedDataIn[500] = 0;
decompressedDataIn[501] = 0;
decompressedDataIn[502] = 0;
decompressedDataIn[503] = 0;
decompressedDataIn[504] = 1;
decompressedDataIn[505] = 0;
decompressedDataIn[506] = 0;
decompressedDataIn[507] = 0;
decompressedDataIn[508] = 0;
decompressedDataIn[509] = 0;
decompressedDataIn[510] = 0;
decompressedDataIn[511] = 0;
decompressedDataIn[512] = 1;
decompressedDataIn[513] = 0;
decompressedDataIn[514] = 0;
decompressedDataIn[515] = 0;
decompressedDataIn[516] = 4;
decompressedDataIn[517] = 0;
decompressedDataIn[518] = 0;
decompressedDataIn[519] = 0;
decompressedDataIn[520] = 4;
decompressedDataIn[521] = 114;
decompressedDataIn[522] = 218;
decompressedDataIn[523] = 23;
decompressedDataIn[524] = 0;
decompressedDataIn[525] = 0;
decompressedDataIn[526] = 0;
decompressedDataIn[527] = 0;
decompressedDataIn[528] = 0;
decompressedDataIn[529] = 224;
decompressedDataIn[530] = 87;
decompressedDataIn[531] = 247;
decompressedDataIn[532] = 217;
decompressedDataIn[533] = 127;
decompressedDataIn[534] = 0;
decompressedDataIn[535] = 0;
decompressedDataIn[536] = 0;
decompressedDataIn[537] = 0;
decompressedDataIn[538] = 0;
decompressedDataIn[539] = 0;
decompressedDataIn[540] = 0;
decompressedDataIn[541] = 0;
decompressedDataIn[542] = 0;
decompressedDataIn[543] = 0;
decompressedDataIn[544] = 0;
decompressedDataIn[545] = 16;
decompressedDataIn[546] = 0;
decompressedDataIn[547] = 0;
decompressedDataIn[548] = 0;
decompressedDataIn[549] = 0;
decompressedDataIn[550] = 0;
decompressedDataIn[551] = 0;
decompressedDataIn[552] = 0;
decompressedDataIn[553] = 16;
decompressedDataIn[554] = 0;
decompressedDataIn[555] = 0;
decompressedDataIn[556] = 0;
decompressedDataIn[557] = 0;
decompressedDataIn[558] = 0;
decompressedDataIn[559] = 0;
decompressedDataIn[560] = 1;
decompressedDataIn[561] = 0;
decompressedDataIn[562] = 0;
decompressedDataIn[563] = 0;
decompressedDataIn[564] = 0;
decompressedDataIn[565] = 0;
decompressedDataIn[566] = 0;
decompressedDataIn[567] = 0;
decompressedDataIn[568] = 1;
decompressedDataIn[569] = 0;
decompressedDataIn[570] = 0;
decompressedDataIn[571] = 0;
decompressedDataIn[572] = 6;
decompressedDataIn[573] = 0;
decompressedDataIn[574] = 0;
decompressedDataIn[575] = 0;
decompressedDataIn[576] = 4;
decompressedDataIn[577] = 130;
decompressedDataIn[578] = 218;
decompressedDataIn[579] = 23;
decompressedDataIn[580] = 0;
decompressedDataIn[581] = 0;
decompressedDataIn[582] = 0;
decompressedDataIn[583] = 0;
decompressedDataIn[584] = 0;
decompressedDataIn[585] = 240;
decompressedDataIn[586] = 87;
decompressedDataIn[587] = 247;
decompressedDataIn[588] = 217;
decompressedDataIn[589] = 127;
decompressedDataIn[590] = 0;
decompressedDataIn[591] = 0;
decompressedDataIn[592] = 0;
decompressedDataIn[593] = 0;
decompressedDataIn[594] = 0;
decompressedDataIn[595] = 0;
decompressedDataIn[596] = 0;
decompressedDataIn[597] = 0;
decompressedDataIn[598] = 0;
decompressedDataIn[599] = 0;
decompressedDataIn[600] = 0;
decompressedDataIn[601] = 16;
decompressedDataIn[602] = 0;
decompressedDataIn[603] = 0;
decompressedDataIn[604] = 0;
decompressedDataIn[605] = 0;
decompressedDataIn[606] = 0;
decompressedDataIn[607] = 0;
decompressedDataIn[608] = 0;
decompressedDataIn[609] = 16;
decompressedDataIn[610] = 0;
decompressedDataIn[611] = 0;
decompressedDataIn[612] = 0;
decompressedDataIn[613] = 0;
decompressedDataIn[614] = 0;
decompressedDataIn[615] = 0;
decompressedDataIn[616] = 1;
decompressedDataIn[617] = 0;
decompressedDataIn[618] = 0;
decompressedDataIn[619] = 0;
decompressedDataIn[620] = 0;
decompressedDataIn[621] = 0;
decompressedDataIn[622] = 0;
decompressedDataIn[623] = 0;
decompressedDataIn[624] = 1;
decompressedDataIn[625] = 0;
decompressedDataIn[626] = 0;
decompressedDataIn[627] = 0;
decompressedDataIn[628] = 6;
decompressedDataIn[629] = 0;
decompressedDataIn[630] = 0;
decompressedDataIn[631] = 0;
decompressedDataIn[632] = 4;
decompressedDataIn[633] = 146;
decompressedDataIn[634] = 218;
decompressedDataIn[635] = 23;
decompressedDataIn[636] = 0;
decompressedDataIn[637] = 0;
decompressedDataIn[638] = 0;
decompressedDataIn[639] = 0;
decompressedDataIn[640] = 0;
decompressedDataIn[641] = 0;
decompressedDataIn[642] = 88;
decompressedDataIn[643] = 247;
decompressedDataIn[644] = 217;
decompressedDataIn[645] = 127;
decompressedDataIn[646] = 0;
decompressedDataIn[647] = 0;
decompressedDataIn[648] = 0;
decompressedDataIn[649] = 0;
decompressedDataIn[650] = 0;
decompressedDataIn[651] = 0;
decompressedDataIn[652] = 0;
decompressedDataIn[653] = 0;
decompressedDataIn[654] = 0;
decompressedDataIn[655] = 0;
decompressedDataIn[656] = 0;
decompressedDataIn[657] = 64;
decompressedDataIn[658] = 0;
decompressedDataIn[659] = 0;
decompressedDataIn[660] = 0;
decompressedDataIn[661] = 0;
decompressedDataIn[662] = 0;
decompressedDataIn[663] = 0;
decompressedDataIn[664] = 0;
decompressedDataIn[665] = 64;
decompressedDataIn[666] = 0;
decompressedDataIn[667] = 0;
decompressedDataIn[668] = 0;
decompressedDataIn[669] = 0;
decompressedDataIn[670] = 0;
decompressedDataIn[671] = 0;
decompressedDataIn[672] = 1;
decompressedDataIn[673] = 0;
decompressedDataIn[674] = 0;
decompressedDataIn[675] = 0;
decompressedDataIn[676] = 0;
decompressedDataIn[677] = 0;
decompressedDataIn[678] = 0;
decompressedDataIn[679] = 0;
decompressedDataIn[680] = 1;
decompressedDataIn[681] = 0;
decompressedDataIn[682] = 0;
decompressedDataIn[683] = 0;
decompressedDataIn[684] = 4;
decompressedDataIn[685] = 0;
decompressedDataIn[686] = 0;
decompressedDataIn[687] = 0;
decompressedDataIn[688] = 4;
decompressedDataIn[689] = 210;
decompressedDataIn[690] = 218;
decompressedDataIn[691] = 23;
decompressedDataIn[692] = 0;
decompressedDataIn[693] = 0;
decompressedDataIn[694] = 0;
decompressedDataIn[695] = 0;
decompressedDataIn[696] = 0;
decompressedDataIn[697] = 0;
decompressedDataIn[698] = 146;
decompressedDataIn[699] = 247;
decompressedDataIn[700] = 217;
decompressedDataIn[701] = 127;
decompressedDataIn[702] = 0;
decompressedDataIn[703] = 0;
decompressedDataIn[704] = 0;
decompressedDataIn[705] = 0;
decompressedDataIn[706] = 0;
decompressedDataIn[707] = 0;
decompressedDataIn[708] = 0;
decompressedDataIn[709] = 0;
decompressedDataIn[710] = 0;
decompressedDataIn[711] = 0;
decompressedDataIn[712] = 0;
decompressedDataIn[713] = 16;
decompressedDataIn[714] = 0;
decompressedDataIn[715] = 0;
decompressedDataIn[716] = 0;
decompressedDataIn[717] = 0;
decompressedDataIn[718] = 0;
decompressedDataIn[719] = 0;
decompressedDataIn[720] = 0;
decompressedDataIn[721] = 16;
decompressedDataIn[722] = 0;
decompressedDataIn[723] = 0;
decompressedDataIn[724] = 0;
decompressedDataIn[725] = 0;
decompressedDataIn[726] = 0;
decompressedDataIn[727] = 0;
decompressedDataIn[728] = 1;
decompressedDataIn[729] = 0;
decompressedDataIn[730] = 0;
decompressedDataIn[731] = 0;
decompressedDataIn[732] = 0;
decompressedDataIn[733] = 0;
decompressedDataIn[734] = 0;
decompressedDataIn[735] = 0;
decompressedDataIn[736] = 1;
decompressedDataIn[737] = 0;
decompressedDataIn[738] = 0;
decompressedDataIn[739] = 0;
decompressedDataIn[740] = 6;
decompressedDataIn[741] = 0;
decompressedDataIn[742] = 0;
decompressedDataIn[743] = 0;
decompressedDataIn[744] = 4;
decompressedDataIn[745] = 226;
decompressedDataIn[746] = 218;
decompressedDataIn[747] = 23;
decompressedDataIn[748] = 0;
decompressedDataIn[749] = 0;
decompressedDataIn[750] = 0;
decompressedDataIn[751] = 0;
decompressedDataIn[752] = 0;
decompressedDataIn[753] = 16;
decompressedDataIn[754] = 146;
decompressedDataIn[755] = 247;
decompressedDataIn[756] = 217;
decompressedDataIn[757] = 127;
decompressedDataIn[758] = 0;
decompressedDataIn[759] = 0;
decompressedDataIn[760] = 0;
decompressedDataIn[761] = 0;
decompressedDataIn[762] = 0;
decompressedDataIn[763] = 0;
decompressedDataIn[764] = 0;
decompressedDataIn[765] = 0;
decompressedDataIn[766] = 0;
decompressedDataIn[767] = 0;
decompressedDataIn[768] = 0;
decompressedDataIn[769] = 16;
decompressedDataIn[770] = 0;
decompressedDataIn[771] = 0;
decompressedDataIn[772] = 0;
decompressedDataIn[773] = 0;
decompressedDataIn[774] = 0;
decompressedDataIn[775] = 0;
decompressedDataIn[776] = 0;
decompressedDataIn[777] = 16;
decompressedDataIn[778] = 0;
decompressedDataIn[779] = 0;
decompressedDataIn[780] = 0;
decompressedDataIn[781] = 0;
decompressedDataIn[782] = 0;
decompressedDataIn[783] = 0;
decompressedDataIn[784] = 1;
decompressedDataIn[785] = 0;
decompressedDataIn[786] = 0;
decompressedDataIn[787] = 0;
decompressedDataIn[788] = 0;
decompressedDataIn[789] = 0;
decompressedDataIn[790] = 0;
decompressedDataIn[791] = 0;
decompressedDataIn[792] = 1;
decompressedDataIn[793] = 0;
decompressedDataIn[794] = 0;
decompressedDataIn[795] = 0;
decompressedDataIn[796] = 6;
decompressedDataIn[797] = 0;
decompressedDataIn[798] = 0;
decompressedDataIn[799] = 0;
decompressedDataIn[800] = 4;
decompressedDataIn[801] = 242;
decompressedDataIn[802] = 218;
decompressedDataIn[803] = 23;
decompressedDataIn[804] = 0;
decompressedDataIn[805] = 0;
decompressedDataIn[806] = 0;
decompressedDataIn[807] = 0;
decompressedDataIn[808] = 0;
decompressedDataIn[809] = 224;
decompressedDataIn[810] = 178;
decompressedDataIn[811] = 247;
decompressedDataIn[812] = 217;
decompressedDataIn[813] = 127;
decompressedDataIn[814] = 0;
decompressedDataIn[815] = 0;
decompressedDataIn[816] = 0;
decompressedDataIn[817] = 0;
decompressedDataIn[818] = 0;
decompressedDataIn[819] = 0;
decompressedDataIn[820] = 0;
decompressedDataIn[821] = 0;
decompressedDataIn[822] = 0;
decompressedDataIn[823] = 0;
decompressedDataIn[824] = 0;
decompressedDataIn[825] = 80;
decompressedDataIn[826] = 0;
decompressedDataIn[827] = 0;
decompressedDataIn[828] = 0;
decompressedDataIn[829] = 0;
decompressedDataIn[830] = 0;
decompressedDataIn[831] = 0;
decompressedDataIn[832] = 0;
decompressedDataIn[833] = 80;
decompressedDataIn[834] = 0;
decompressedDataIn[835] = 0;
decompressedDataIn[836] = 0;
decompressedDataIn[837] = 0;
decompressedDataIn[838] = 0;
decompressedDataIn[839] = 0;
decompressedDataIn[840] = 1;
decompressedDataIn[841] = 0;
decompressedDataIn[842] = 0;
decompressedDataIn[843] = 0;
decompressedDataIn[844] = 0;
decompressedDataIn[845] = 0;
decompressedDataIn[846] = 0;
decompressedDataIn[847] = 0;
decompressedDataIn[848] = 1;
decompressedDataIn[849] = 0;
decompressedDataIn[850] = 0;
decompressedDataIn[851] = 0;
decompressedDataIn[852] = 4;
decompressedDataIn[853] = 0;
decompressedDataIn[854] = 0;
decompressedDataIn[855] = 0;
decompressedDataIn[856] = 4;
decompressedDataIn[857] = 66;
decompressedDataIn[858] = 219;
decompressedDataIn[859] = 23;
decompressedDataIn[860] = 0;
decompressedDataIn[861] = 0;
decompressedDataIn[862] = 0;
decompressedDataIn[863] = 0;
decompressedDataIn[864] = 0;
decompressedDataIn[865] = 144;
decompressedDataIn[866] = 180;
decompressedDataIn[867] = 247;
decompressedDataIn[868] = 217;
decompressedDataIn[869] = 127;
decompressedDataIn[870] = 0;
decompressedDataIn[871] = 0;
decompressedDataIn[872] = 0;
decompressedDataIn[873] = 0;
decompressedDataIn[874] = 0;
decompressedDataIn[875] = 0;
decompressedDataIn[876] = 0;
decompressedDataIn[877] = 0;
decompressedDataIn[878] = 0;
decompressedDataIn[879] = 0;
decompressedDataIn[880] = 0;
decompressedDataIn[881] = 16;
decompressedDataIn[882] = 0;
decompressedDataIn[883] = 0;
decompressedDataIn[884] = 0;
decompressedDataIn[885] = 0;
decompressedDataIn[886] = 0;
decompressedDataIn[887] = 0;
decompressedDataIn[888] = 0;
decompressedDataIn[889] = 16;
decompressedDataIn[890] = 0;
decompressedDataIn[891] = 0;
decompressedDataIn[892] = 0;
decompressedDataIn[893] = 0;
decompressedDataIn[894] = 0;
decompressedDataIn[895] = 0;
decompressedDataIn[896] = 1;
decompressedDataIn[897] = 0;
decompressedDataIn[898] = 0;
decompressedDataIn[899] = 0;
decompressedDataIn[900] = 0;
decompressedDataIn[901] = 0;
decompressedDataIn[902] = 0;
decompressedDataIn[903] = 0;
decompressedDataIn[904] = 1;
decompressedDataIn[905] = 0;
decompressedDataIn[906] = 0;
decompressedDataIn[907] = 0;
decompressedDataIn[908] = 6;
decompressedDataIn[909] = 0;
decompressedDataIn[910] = 0;
decompressedDataIn[911] = 0;
decompressedDataIn[912] = 4;
decompressedDataIn[913] = 82;
decompressedDataIn[914] = 219;
decompressedDataIn[915] = 23;
decompressedDataIn[916] = 0;
decompressedDataIn[917] = 0;
decompressedDataIn[918] = 0;
decompressedDataIn[919] = 0;
decompressedDataIn[920] = 0;
decompressedDataIn[921] = 160;
decompressedDataIn[922] = 180;
decompressedDataIn[923] = 247;
decompressedDataIn[924] = 217;
decompressedDataIn[925] = 127;
decompressedDataIn[926] = 0;
decompressedDataIn[927] = 0;
decompressedDataIn[928] = 0;
decompressedDataIn[929] = 0;
decompressedDataIn[930] = 0;
decompressedDataIn[931] = 0;
decompressedDataIn[932] = 0;
decompressedDataIn[933] = 0;
decompressedDataIn[934] = 0;
decompressedDataIn[935] = 0;
decompressedDataIn[936] = 0;
decompressedDataIn[937] = 16;
decompressedDataIn[938] = 0;
decompressedDataIn[939] = 0;
decompressedDataIn[940] = 0;
decompressedDataIn[941] = 0;
decompressedDataIn[942] = 0;
decompressedDataIn[943] = 0;
decompressedDataIn[944] = 0;
decompressedDataIn[945] = 16;
decompressedDataIn[946] = 0;
decompressedDataIn[947] = 0;
decompressedDataIn[948] = 0;
decompressedDataIn[949] = 0;
decompressedDataIn[950] = 0;
decompressedDataIn[951] = 0;
decompressedDataIn[952] = 1;
decompressedDataIn[953] = 0;
decompressedDataIn[954] = 0;
decompressedDataIn[955] = 0;
decompressedDataIn[956] = 0;
decompressedDataIn[957] = 0;
decompressedDataIn[958] = 0;
decompressedDataIn[959] = 0;
decompressedDataIn[960] = 1;
decompressedDataIn[961] = 0;
decompressedDataIn[962] = 0;
decompressedDataIn[963] = 0;
decompressedDataIn[964] = 6;
decompressedDataIn[965] = 0;
decompressedDataIn[966] = 0;
decompressedDataIn[967] = 0;
decompressedDataIn[968] = 4;
decompressedDataIn[969] = 98;
decompressedDataIn[970] = 219;
decompressedDataIn[971] = 23;
decompressedDataIn[972] = 0;
decompressedDataIn[973] = 0;
decompressedDataIn[974] = 0;
decompressedDataIn[975] = 0;
decompressedDataIn[976] = 0;
decompressedDataIn[977] = 176;
decompressedDataIn[978] = 180;
decompressedDataIn[979] = 247;
decompressedDataIn[980] = 217;
decompressedDataIn[981] = 127;
decompressedDataIn[982] = 0;
decompressedDataIn[983] = 0;
decompressedDataIn[984] = 0;
decompressedDataIn[985] = 0;
decompressedDataIn[986] = 0;
decompressedDataIn[987] = 0;
decompressedDataIn[988] = 0;
decompressedDataIn[989] = 0;
decompressedDataIn[990] = 0;
decompressedDataIn[991] = 0;
decompressedDataIn[992] = 0;
decompressedDataIn[993] = 16;
decompressedDataIn[994] = 0;
decompressedDataIn[995] = 0;
decompressedDataIn[996] = 0;
decompressedDataIn[997] = 0;
decompressedDataIn[998] = 0;
decompressedDataIn[999] = 0;
decompressedDataIn[1000] = 0;
decompressedDataIn[1001] = 16;
decompressedDataIn[1002] = 0;
decompressedDataIn[1003] = 0;
decompressedDataIn[1004] = 0;
decompressedDataIn[1005] = 0;
decompressedDataIn[1006] = 0;
decompressedDataIn[1007] = 0;
decompressedDataIn[1008] = 1;
decompressedDataIn[1009] = 0;
decompressedDataIn[1010] = 0;
decompressedDataIn[1011] = 0;
decompressedDataIn[1012] = 0;
decompressedDataIn[1013] = 0;
decompressedDataIn[1014] = 0;
decompressedDataIn[1015] = 0;
decompressedDataIn[1016] = 1;
decompressedDataIn[1017] = 0;
decompressedDataIn[1018] = 0;
decompressedDataIn[1019] = 0;
decompressedDataIn[1020] = 6;
decompressedDataIn[1021] = 0;
decompressedDataIn[1022] = 0;
decompressedDataIn[1023] = 0;
decompressedDataIn[1024] = 4;
decompressedDataIn[1025] = 114;
decompressedDataIn[1026] = 219;
decompressedDataIn[1027] = 23;
decompressedDataIn[1028] = 0;
decompressedDataIn[1029] = 0;
decompressedDataIn[1030] = 0;
decompressedDataIn[1031] = 0;
decompressedDataIn[1032] = 0;
decompressedDataIn[1033] = 128;
decompressedDataIn[1034] = 65;
decompressedDataIn[1035] = 67;
decompressedDataIn[1036] = 255;
decompressedDataIn[1037] = 127;
decompressedDataIn[1038] = 0;
decompressedDataIn[1039] = 0;
decompressedDataIn[1040] = 0;
decompressedDataIn[1041] = 0;
decompressedDataIn[1042] = 0;
decompressedDataIn[1043] = 0;
decompressedDataIn[1044] = 0;
decompressedDataIn[1045] = 0;
decompressedDataIn[1046] = 0;
decompressedDataIn[1047] = 0;
decompressedDataIn[1048] = 0;
decompressedDataIn[1049] = 16;
decompressedDataIn[1050] = 2;
decompressedDataIn[1051] = 0;
decompressedDataIn[1052] = 0;
decompressedDataIn[1053] = 0;
decompressedDataIn[1054] = 0;
decompressedDataIn[1055] = 0;
decompressedDataIn[1056] = 0;
decompressedDataIn[1057] = 16;
decompressedDataIn[1058] = 2;
decompressedDataIn[1059] = 0;
decompressedDataIn[1060] = 0;
decompressedDataIn[1061] = 0;
decompressedDataIn[1062] = 0;
decompressedDataIn[1063] = 0;
decompressedDataIn[1064] = 1;
decompressedDataIn[1065] = 0;
decompressedDataIn[1066] = 0;
decompressedDataIn[1067] = 0;
decompressedDataIn[1068] = 0;
decompressedDataIn[1069] = 0;
decompressedDataIn[1070] = 0;
decompressedDataIn[1071] = 0;
decompressedDataIn[1072] = 1;
decompressedDataIn[1073] = 0;
decompressedDataIn[1074] = 0;
decompressedDataIn[1075] = 0;
decompressedDataIn[1076] = 5;
decompressedDataIn[1077] = 0;
decompressedDataIn[1078] = 0;
decompressedDataIn[1079] = 0;
decompressedDataIn[1080] = 4;
decompressedDataIn[1081] = 130;
decompressedDataIn[1082] = 221;
decompressedDataIn[1083] = 23;
decompressedDataIn[1084] = 0;
decompressedDataIn[1085] = 0;
decompressedDataIn[1086] = 0;
decompressedDataIn[1087] = 0;
decompressedDataIn[1088] = 0;
decompressedDataIn[1089] = 64;
decompressedDataIn[1090] = 94;
decompressedDataIn[1091] = 67;
decompressedDataIn[1092] = 255;
decompressedDataIn[1093] = 127;
decompressedDataIn[1094] = 0;
decompressedDataIn[1095] = 0;
decompressedDataIn[1096] = 0;
decompressedDataIn[1097] = 0;
decompressedDataIn[1098] = 0;
decompressedDataIn[1099] = 0;
decompressedDataIn[1100] = 0;
decompressedDataIn[1101] = 0;
decompressedDataIn[1102] = 0;
decompressedDataIn[1103] = 0;
decompressedDataIn[1104] = 0;
decompressedDataIn[1105] = 16;
decompressedDataIn[1106] = 0;
decompressedDataIn[1107] = 0;
decompressedDataIn[1108] = 0;
decompressedDataIn[1109] = 0;
decompressedDataIn[1110] = 0;
decompressedDataIn[1111] = 0;
decompressedDataIn[1112] = 0;
decompressedDataIn[1113] = 16;
decompressedDataIn[1114] = 0;
decompressedDataIn[1115] = 0;
decompressedDataIn[1116] = 0;
decompressedDataIn[1117] = 0;
decompressedDataIn[1118] = 0;
decompressedDataIn[1119] = 0;
decompressedDataIn[1120] = 1;
decompressedDataIn[1121] = 0;
decompressedDataIn[1122] = 0;
decompressedDataIn[1123] = 0;
decompressedDataIn[1124] = 0;
decompressedDataIn[1125] = 0;
decompressedDataIn[1126] = 0;
decompressedDataIn[1127] = 0;
decompressedDataIn[1128] = 1;
decompressedDataIn[1129] = 0;
decompressedDataIn[1130] = 0;
decompressedDataIn[1131] = 0;
decompressedDataIn[1132] = 5;
decompressedDataIn[1133] = 0;
decompressedDataIn[1134] = 0;
decompressedDataIn[1135] = 0;
decompressedDataIn[1136] = 4;
decompressedDataIn[1137] = 146;
decompressedDataIn[1138] = 221;
decompressedDataIn[1139] = 23;
decompressedDataIn[1140] = 0;
decompressedDataIn[1141] = 0;
decompressedDataIn[1142] = 0;
decompressedDataIn[1143] = 0;
decompressedDataIn[1144] = 0;
decompressedDataIn[1145] = 0;
decompressedDataIn[1146] = 96;
decompressedDataIn[1147] = 255;
decompressedDataIn[1148] = 255;
decompressedDataIn[1149] = 255;
decompressedDataIn[1150] = 255;
decompressedDataIn[1151] = 255;
decompressedDataIn[1152] = 0;
decompressedDataIn[1153] = 0;
decompressedDataIn[1154] = 0;
decompressedDataIn[1155] = 0;
decompressedDataIn[1156] = 0;
decompressedDataIn[1157] = 0;
decompressedDataIn[1158] = 0;
decompressedDataIn[1159] = 0;
decompressedDataIn[1160] = 0;
decompressedDataIn[1161] = 16;
decompressedDataIn[1162] = 0;
decompressedDataIn[1163] = 0;
decompressedDataIn[1164] = 0;
decompressedDataIn[1165] = 0;
decompressedDataIn[1166] = 0;
decompressedDataIn[1167] = 0;
decompressedDataIn[1168] = 0;
decompressedDataIn[1169] = 16;
decompressedDataIn[1170] = 0;
decompressedDataIn[1171] = 0;
decompressedDataIn[1172] = 0;
decompressedDataIn[1173] = 0;
decompressedDataIn[1174] = 0;
decompressedDataIn[1175] = 0;
decompressedDataIn[1176] = 1;
decompressedDataIn[1177] = 0;
decompressedDataIn[1178] = 0;
decompressedDataIn[1179] = 0;
decompressedDataIn[1180] = 0;
decompressedDataIn[1181] = 0;
decompressedDataIn[1182] = 0;
decompressedDataIn[1183] = 0;
decompressedDataIn[1184] = 5;
decompressedDataIn[1185] = 0;
decompressedDataIn[1186] = 0;
decompressedDataIn[1187] = 0;
decompressedDataIn[1188] = 136;
decompressedDataIn[1189] = 0;
decompressedDataIn[1190] = 0;
decompressedDataIn[1191] = 0;
decompressedDataIn[1192] = 3;
decompressedDataIn[1193] = 0;
decompressedDataIn[1194] = 0;
decompressedDataIn[1195] = 0;
decompressedDataIn[1196] = 67;
decompressedDataIn[1197] = 79;
decompressedDataIn[1198] = 82;
decompressedDataIn[1199] = 69;
decompressedDataIn[1200] = 0;
decompressedDataIn[1201] = 0;
decompressedDataIn[1202] = 0;
decompressedDataIn[1203] = 0;
decompressedDataIn[1204] = 0;
decompressedDataIn[1205] = 116;
decompressedDataIn[1206] = 0;
decompressedDataIn[1207] = 0;
decompressedDataIn[1208] = 0;
decompressedDataIn[1209] = 0;
decompressedDataIn[1210] = 0;
decompressedDataIn[1211] = 0;
decompressedDataIn[1212] = 0;
decompressedDataIn[1213] = 0;
decompressedDataIn[1214] = 64;
decompressedDataIn[1215] = 64;
decompressedDataIn[1216] = 0;
decompressedDataIn[1217] = 0;
decompressedDataIn[1218] = 0;
decompressedDataIn[1219] = 0;
decompressedDataIn[1220] = 0;
decompressedDataIn[1221] = 0;
decompressedDataIn[1222] = 0;
decompressedDataIn[1223] = 0;
decompressedDataIn[1224] = 0;
decompressedDataIn[1225] = 0;
decompressedDataIn[1226] = 0;
decompressedDataIn[1227] = 0;
decompressedDataIn[1228] = 237;
decompressedDataIn[1229] = 17;
decompressedDataIn[1230] = 0;
decompressedDataIn[1231] = 0;
decompressedDataIn[1232] = 234;
decompressedDataIn[1233] = 17;
decompressedDataIn[1234] = 0;
decompressedDataIn[1235] = 0;
decompressedDataIn[1236] = 147;
decompressedDataIn[1237] = 16;
decompressedDataIn[1238] = 0;
decompressedDataIn[1239] = 0;
decompressedDataIn[1240] = 116;
decompressedDataIn[1241] = 12;
decompressedDataIn[1242] = 0;
decompressedDataIn[1243] = 0;
decompressedDataIn[1244] = 98;
decompressedDataIn[1245] = 108;
decompressedDataIn[1246] = 97;
decompressedDataIn[1247] = 99;
decompressedDataIn[1248] = 107;
decompressedDataIn[1249] = 115;
decompressedDataIn[1250] = 99;
decompressedDataIn[1251] = 104;
decompressedDataIn[1252] = 111;
decompressedDataIn[1253] = 108;
decompressedDataIn[1254] = 101;
decompressedDataIn[1255] = 115;
decompressedDataIn[1256] = 0;
decompressedDataIn[1257] = 0;
decompressedDataIn[1258] = 0;
decompressedDataIn[1259] = 0;
decompressedDataIn[1260] = 47;
decompressedDataIn[1261] = 104;
decompressedDataIn[1262] = 111;
decompressedDataIn[1263] = 109;
decompressedDataIn[1264] = 101;
decompressedDataIn[1265] = 47;
decompressedDataIn[1266] = 118;
decompressedDataIn[1267] = 116;
decompressedDataIn[1268] = 45;
decompressedDataIn[1269] = 99;
decompressedDataIn[1270] = 115;
decompressedDataIn[1271] = 47;
decompressedDataIn[1272] = 109;
decompressedDataIn[1273] = 108;
decompressedDataIn[1274] = 97;
decompressedDataIn[1275] = 103;
decompressedDataIn[1276] = 104;
decompressedDataIn[1277] = 97;
decompressedDataIn[1278] = 114;
decompressedDataIn[1279] = 105;
decompressedDataIn[1280] = 47;
decompressedDataIn[1281] = 112;
decompressedDataIn[1282] = 97;
decompressedDataIn[1283] = 114;
decompressedDataIn[1284] = 115;
decompressedDataIn[1285] = 101;
decompressedDataIn[1286] = 99;
decompressedDataIn[1287] = 45;
decompressedDataIn[1288] = 98;
decompressedDataIn[1289] = 101;
decompressedDataIn[1290] = 110;
decompressedDataIn[1291] = 99;
decompressedDataIn[1292] = 104;
decompressedDataIn[1293] = 109;
decompressedDataIn[1294] = 97;
decompressedDataIn[1295] = 114;
decompressedDataIn[1296] = 107;
decompressedDataIn[1297] = 95;
decompressedDataIn[1298] = 110;
decompressedDataIn[1299] = 118;
decompressedDataIn[1300] = 109;
decompressedDataIn[1301] = 101;
decompressedDataIn[1302] = 95;
decompressedDataIn[1303] = 114;
decompressedDataIn[1304] = 101;
decompressedDataIn[1305] = 115;
decompressedDataIn[1306] = 117;
decompressedDataIn[1307] = 108;
decompressedDataIn[1308] = 116;
decompressedDataIn[1309] = 115;
decompressedDataIn[1310] = 47;
decompressedDataIn[1311] = 112;
decompressedDataIn[1312] = 107;
decompressedDataIn[1313] = 103;
decompressedDataIn[1314] = 115;
decompressedDataIn[1315] = 47;
decompressedDataIn[1316] = 97;
decompressedDataIn[1317] = 112;
decompressedDataIn[1318] = 112;
decompressedDataIn[1319] = 115;
decompressedDataIn[1320] = 47;
decompressedDataIn[1321] = 98;
decompressedDataIn[1322] = 108;
decompressedDataIn[1323] = 97;
decompressedDataIn[1324] = 99;
decompressedDataIn[1325] = 107;
decompressedDataIn[1326] = 115;
decompressedDataIn[1327] = 99;
decompressedDataIn[1328] = 104;
decompressedDataIn[1329] = 111;
decompressedDataIn[1330] = 108;
decompressedDataIn[1331] = 101;
decompressedDataIn[1332] = 115;
decompressedDataIn[1333] = 47;
decompressedDataIn[1334] = 105;
decompressedDataIn[1335] = 110;
decompressedDataIn[1336] = 115;
decompressedDataIn[1337] = 116;
decompressedDataIn[1338] = 47;
decompressedDataIn[1339] = 97;
decompressedDataIn[1340] = 5;
decompressedDataIn[1341] = 0;
decompressedDataIn[1342] = 0;
decompressedDataIn[1343] = 0;
decompressedDataIn[1344] = 80;
decompressedDataIn[1345] = 1;
decompressedDataIn[1346] = 0;
decompressedDataIn[1347] = 0;
decompressedDataIn[1348] = 1;
decompressedDataIn[1349] = 0;
decompressedDataIn[1350] = 0;
decompressedDataIn[1351] = 0;
decompressedDataIn[1352] = 67;
decompressedDataIn[1353] = 79;
decompressedDataIn[1354] = 82;
decompressedDataIn[1355] = 69;
decompressedDataIn[1356] = 0;
decompressedDataIn[1357] = 0;
decompressedDataIn[1358] = 0;
decompressedDataIn[1359] = 0;
decompressedDataIn[1360] = 0;
decompressedDataIn[1361] = 0;
decompressedDataIn[1362] = 0;
decompressedDataIn[1363] = 0;
decompressedDataIn[1364] = 0;
decompressedDataIn[1365] = 0;
decompressedDataIn[1366] = 0;
decompressedDataIn[1367] = 0;
decompressedDataIn[1368] = 0;
decompressedDataIn[1369] = 0;
decompressedDataIn[1370] = 0;
decompressedDataIn[1371] = 0;
decompressedDataIn[1372] = 0;
decompressedDataIn[1373] = 0;
decompressedDataIn[1374] = 0;
decompressedDataIn[1375] = 0;
decompressedDataIn[1376] = 0;
decompressedDataIn[1377] = 0;
decompressedDataIn[1378] = 0;
decompressedDataIn[1379] = 0;
decompressedDataIn[1380] = 0;
decompressedDataIn[1381] = 0;
decompressedDataIn[1382] = 0;
decompressedDataIn[1383] = 0;
decompressedDataIn[1384] = 0;
decompressedDataIn[1385] = 0;
decompressedDataIn[1386] = 0;
decompressedDataIn[1387] = 0;
decompressedDataIn[1388] = 0;
decompressedDataIn[1389] = 0;
decompressedDataIn[1390] = 0;
decompressedDataIn[1391] = 0;
decompressedDataIn[1392] = 237;
decompressedDataIn[1393] = 17;
decompressedDataIn[1394] = 0;
decompressedDataIn[1395] = 0;
decompressedDataIn[1396] = 0;
decompressedDataIn[1397] = 0;
decompressedDataIn[1398] = 0;
decompressedDataIn[1399] = 0;
decompressedDataIn[1400] = 0;
decompressedDataIn[1401] = 0;
decompressedDataIn[1402] = 0;
decompressedDataIn[1403] = 0;
decompressedDataIn[1404] = 0;
decompressedDataIn[1405] = 0;
decompressedDataIn[1406] = 0;
decompressedDataIn[1407] = 0;
decompressedDataIn[1408] = 0;
decompressedDataIn[1409] = 0;
decompressedDataIn[1410] = 0;
decompressedDataIn[1411] = 0;
decompressedDataIn[1412] = 0;
decompressedDataIn[1413] = 0;
decompressedDataIn[1414] = 0;
decompressedDataIn[1415] = 0;
decompressedDataIn[1416] = 0;
decompressedDataIn[1417] = 0;
decompressedDataIn[1418] = 0;
decompressedDataIn[1419] = 0;
decompressedDataIn[1420] = 0;
decompressedDataIn[1421] = 0;
decompressedDataIn[1422] = 0;
decompressedDataIn[1423] = 0;
decompressedDataIn[1424] = 0;
decompressedDataIn[1425] = 0;
decompressedDataIn[1426] = 0;
decompressedDataIn[1427] = 0;
decompressedDataIn[1428] = 0;
decompressedDataIn[1429] = 0;
decompressedDataIn[1430] = 0;
decompressedDataIn[1431] = 0;
decompressedDataIn[1432] = 0;
decompressedDataIn[1433] = 0;
decompressedDataIn[1434] = 0;
decompressedDataIn[1435] = 0;
decompressedDataIn[1436] = 0;
decompressedDataIn[1437] = 0;
decompressedDataIn[1438] = 0;
decompressedDataIn[1439] = 0;
decompressedDataIn[1440] = 0;
decompressedDataIn[1441] = 0;
decompressedDataIn[1442] = 0;
decompressedDataIn[1443] = 0;
decompressedDataIn[1444] = 0;
decompressedDataIn[1445] = 0;
decompressedDataIn[1446] = 0;
decompressedDataIn[1447] = 0;
decompressedDataIn[1448] = 0;
decompressedDataIn[1449] = 0;
decompressedDataIn[1450] = 0;
decompressedDataIn[1451] = 0;
decompressedDataIn[1452] = 0;
decompressedDataIn[1453] = 0;
decompressedDataIn[1454] = 0;
decompressedDataIn[1455] = 0;
decompressedDataIn[1456] = 0;
decompressedDataIn[1457] = 0;
decompressedDataIn[1458] = 0;
decompressedDataIn[1459] = 0;
decompressedDataIn[1460] = 0;
decompressedDataIn[1461] = 0;
decompressedDataIn[1462] = 0;
decompressedDataIn[1463] = 0;
decompressedDataIn[1464] = 0;
decompressedDataIn[1465] = 0;
decompressedDataIn[1466] = 0;
decompressedDataIn[1467] = 0;
decompressedDataIn[1468] = 0;
decompressedDataIn[1469] = 0;
decompressedDataIn[1470] = 0;
decompressedDataIn[1471] = 0;
decompressedDataIn[1472] = 1;
decompressedDataIn[1473] = 0;
decompressedDataIn[1474] = 0;
decompressedDataIn[1475] = 0;
decompressedDataIn[1476] = 0;
decompressedDataIn[1477] = 0;
decompressedDataIn[1478] = 0;
decompressedDataIn[1479] = 0;
decompressedDataIn[1480] = 219;
decompressedDataIn[1481] = 177;
decompressedDataIn[1482] = 251;
decompressedDataIn[1483] = 246;
decompressedDataIn[1484] = 217;
decompressedDataIn[1485] = 127;
decompressedDataIn[1486] = 0;
decompressedDataIn[1487] = 0;
decompressedDataIn[1488] = 0;
decompressedDataIn[1489] = 0;
decompressedDataIn[1490] = 0;
decompressedDataIn[1491] = 0;
decompressedDataIn[1492] = 0;
decompressedDataIn[1493] = 0;
decompressedDataIn[1494] = 0;
decompressedDataIn[1495] = 0;
decompressedDataIn[1496] = 1;
decompressedDataIn[1497] = 0;
decompressedDataIn[1498] = 0;
decompressedDataIn[1499] = 0;
decompressedDataIn[1500] = 0;
decompressedDataIn[1501] = 0;
decompressedDataIn[1502] = 0;
decompressedDataIn[1503] = 0;
decompressedDataIn[1504] = 0;
decompressedDataIn[1505] = 0;
decompressedDataIn[1506] = 0;
decompressedDataIn[1507] = 0;
decompressedDataIn[1508] = 0;
decompressedDataIn[1509] = 0;
decompressedDataIn[1510] = 0;
decompressedDataIn[1511] = 80;
decompressedDataIn[1512] = 0;
decompressedDataIn[1513] = 0;
decompressedDataIn[1514] = 0;
decompressedDataIn[1515] = 0;
decompressedDataIn[1516] = 0;
decompressedDataIn[1517] = 0;
decompressedDataIn[1518] = 0;
decompressedDataIn[1519] = 0;
decompressedDataIn[1520] = 255;
decompressedDataIn[1521] = 255;
decompressedDataIn[1522] = 255;
decompressedDataIn[1523] = 255;
decompressedDataIn[1524] = 255;
decompressedDataIn[1525] = 255;
decompressedDataIn[1526] = 255;
decompressedDataIn[1527] = 255;
decompressedDataIn[1528] = 0;
decompressedDataIn[1529] = 0;
decompressedDataIn[1530] = 0;
decompressedDataIn[1531] = 0;
decompressedDataIn[1532] = 0;
decompressedDataIn[1533] = 0;
decompressedDataIn[1534] = 0;
decompressedDataIn[1535] = 0;
decompressedDataIn[1536] = 0;
decompressedDataIn[1537] = 0;
decompressedDataIn[1538] = 0;
decompressedDataIn[1539] = 0;
decompressedDataIn[1540] = 0;
decompressedDataIn[1541] = 0;
decompressedDataIn[1542] = 0;
decompressedDataIn[1543] = 80;
decompressedDataIn[1544] = 0;
decompressedDataIn[1545] = 0;
decompressedDataIn[1546] = 0;
decompressedDataIn[1547] = 0;
decompressedDataIn[1548] = 0;
decompressedDataIn[1549] = 0;
decompressedDataIn[1550] = 0;
decompressedDataIn[1551] = 0;
decompressedDataIn[1552] = 0;
decompressedDataIn[1553] = 0;
decompressedDataIn[1554] = 0;
decompressedDataIn[1555] = 0;
decompressedDataIn[1556] = 0;
decompressedDataIn[1557] = 0;
decompressedDataIn[1558] = 0;
decompressedDataIn[1559] = 128;
decompressedDataIn[1560] = 64;
decompressedDataIn[1561] = 0;
decompressedDataIn[1562] = 0;
decompressedDataIn[1563] = 0;
decompressedDataIn[1564] = 0;
decompressedDataIn[1565] = 0;
decompressedDataIn[1566] = 0;
decompressedDataIn[1567] = 0;
decompressedDataIn[1568] = 0;
decompressedDataIn[1569] = 0;
decompressedDataIn[1570] = 0;
decompressedDataIn[1571] = 0;
decompressedDataIn[1572] = 0;
decompressedDataIn[1573] = 0;
decompressedDataIn[1574] = 0;
decompressedDataIn[1575] = 0;
decompressedDataIn[1576] = 0;
decompressedDataIn[1577] = 0;
decompressedDataIn[1578] = 0;
decompressedDataIn[1579] = 0;
decompressedDataIn[1580] = 0;
decompressedDataIn[1581] = 0;
decompressedDataIn[1582] = 0;
decompressedDataIn[1583] = 160;
decompressedDataIn[1584] = 0;
decompressedDataIn[1585] = 0;
decompressedDataIn[1586] = 0;
decompressedDataIn[1587] = 0;
decompressedDataIn[1588] = 0;
decompressedDataIn[1589] = 0;
decompressedDataIn[1590] = 0;
decompressedDataIn[1591] = 0;
decompressedDataIn[1592] = 2;
decompressedDataIn[1593] = 255;
decompressedDataIn[1594] = 255;
decompressedDataIn[1595] = 255;
decompressedDataIn[1596] = 255;
decompressedDataIn[1597] = 255;
decompressedDataIn[1598] = 255;
decompressedDataIn[1599] = 255;
decompressedDataIn[1600] = 110;
decompressedDataIn[1601] = 196;
decompressedDataIn[1602] = 251;
decompressedDataIn[1603] = 246;
decompressedDataIn[1604] = 217;
decompressedDataIn[1605] = 127;
decompressedDataIn[1606] = 0;
decompressedDataIn[1607] = 0;
decompressedDataIn[1608] = 51;
decompressedDataIn[1609] = 0;
decompressedDataIn[1610] = 0;
decompressedDataIn[1611] = 0;
decompressedDataIn[1612] = 225;
decompressedDataIn[1613] = 85;
decompressedDataIn[1614] = 0;
decompressedDataIn[1615] = 0;
decompressedDataIn[1616] = 70;
decompressedDataIn[1617] = 2;
decompressedDataIn[1618] = 0;
decompressedDataIn[1619] = 0;
decompressedDataIn[1620] = 225;
decompressedDataIn[1621] = 85;
decompressedDataIn[1622] = 0;
decompressedDataIn[1623] = 0;
decompressedDataIn[1624] = 192;
decompressedDataIn[1625] = 103;
decompressedDataIn[1626] = 67;
decompressedDataIn[1627] = 67;
decompressedDataIn[1628] = 255;
decompressedDataIn[1629] = 127;
decompressedDataIn[1630] = 0;
decompressedDataIn[1631] = 0;
decompressedDataIn[1632] = 43;
decompressedDataIn[1633] = 0;
decompressedDataIn[1634] = 0;
decompressedDataIn[1635] = 0;
decompressedDataIn[1636] = 225;
decompressedDataIn[1637] = 85;
decompressedDataIn[1638] = 0;
decompressedDataIn[1639] = 0;
decompressedDataIn[1640] = 64;
decompressedDataIn[1641] = 231;
decompressedDataIn[1642] = 178;
decompressedDataIn[1643] = 247;
decompressedDataIn[1644] = 217;
decompressedDataIn[1645] = 127;
decompressedDataIn[1646] = 0;
decompressedDataIn[1647] = 0;
decompressedDataIn[1648] = 0;
decompressedDataIn[1649] = 0;
decompressedDataIn[1650] = 0;
decompressedDataIn[1651] = 0;
decompressedDataIn[1652] = 0;
decompressedDataIn[1653] = 0;
decompressedDataIn[1654] = 0;
decompressedDataIn[1655] = 0;
decompressedDataIn[1656] = 0;
decompressedDataIn[1657] = 0;
decompressedDataIn[1658] = 0;
decompressedDataIn[1659] = 0;
decompressedDataIn[1660] = 225;
decompressedDataIn[1661] = 85;
decompressedDataIn[1662] = 0;
decompressedDataIn[1663] = 0;
decompressedDataIn[1664] = 0;
decompressedDataIn[1665] = 0;
decompressedDataIn[1666] = 0;
decompressedDataIn[1667] = 0;
decompressedDataIn[1668] = 225;
decompressedDataIn[1669] = 85;
decompressedDataIn[1670] = 0;
decompressedDataIn[1671] = 0;
decompressedDataIn[1672] = 0;
decompressedDataIn[1673] = 0;
decompressedDataIn[1674] = 0;
decompressedDataIn[1675] = 0;
decompressedDataIn[1676] = 225;
decompressedDataIn[1677] = 85;
decompressedDataIn[1678] = 0;
decompressedDataIn[1679] = 0;
decompressedDataIn[1680] = 0;
decompressedDataIn[1681] = 0;
decompressedDataIn[1682] = 0;
decompressedDataIn[1683] = 0;
decompressedDataIn[1684] = 225;
decompressedDataIn[1685] = 85;
decompressedDataIn[1686] = 0;
decompressedDataIn[1687] = 0;
decompressedDataIn[1688] = 0;
decompressedDataIn[1689] = 0;
decompressedDataIn[1690] = 0;
decompressedDataIn[1691] = 0;
decompressedDataIn[1692] = 0;
decompressedDataIn[1693] = 0;
decompressedDataIn[1694] = 0;
decompressedDataIn[1695] = 0;
decompressedDataIn[1696] = 5;
decompressedDataIn[1697] = 0;
decompressedDataIn[1698] = 0;
decompressedDataIn[1699] = 0;
decompressedDataIn[1700] = 0;
decompressedDataIn[1701] = 2;
decompressedDataIn[1702] = 0;
decompressedDataIn[1703] = 0;
decompressedDataIn[1704] = 2;
decompressedDataIn[1705] = 0;
decompressedDataIn[1706] = 0;
decompressedDataIn[1707] = 0;
decompressedDataIn[1708] = 67;
decompressedDataIn[1709] = 79;
decompressedDataIn[1710] = 82;
decompressedDataIn[1711] = 69;
decompressedDataIn[1712] = 0;
decompressedDataIn[1713] = 0;
decompressedDataIn[1714] = 0;
decompressedDataIn[1715] = 0;
decompressedDataIn[1716] = 255;
decompressedDataIn[1717] = 255;
decompressedDataIn[1718] = 255;
decompressedDataIn[1719] = 255;
decompressedDataIn[1720] = 255;
decompressedDataIn[1721] = 0;
decompressedDataIn[1722] = 255;
decompressedDataIn[1723] = 7;
decompressedDataIn[1724] = 106;
decompressedDataIn[1725] = 102;
decompressedDataIn[1726] = 14;
decompressedDataIn[1727] = 210;
decompressedDataIn[1728] = 225;
decompressedDataIn[1729] = 85;
decompressedDataIn[1730] = 0;
decompressedDataIn[1731] = 0;
decompressedDataIn[1732] = 0;
decompressedDataIn[1733] = 194;
decompressedDataIn[1734] = 55;
decompressedDataIn[1735] = 75;
decompressedDataIn[1736] = 254;
decompressedDataIn[1737] = 127;
decompressedDataIn[1738] = 0;
decompressedDataIn[1739] = 0;
decompressedDataIn[1740] = 160;
decompressedDataIn[1741] = 31;
decompressedDataIn[1742] = 0;
decompressedDataIn[1743] = 0;
decompressedDataIn[1744] = 0;
decompressedDataIn[1745] = 0;
decompressedDataIn[1746] = 0;
decompressedDataIn[1747] = 0;
decompressedDataIn[1748] = 0;
decompressedDataIn[1749] = 0;
decompressedDataIn[1750] = 0;
decompressedDataIn[1751] = 0;
decompressedDataIn[1752] = 0;
decompressedDataIn[1753] = 0;
decompressedDataIn[1754] = 0;
decompressedDataIn[1755] = 0;
decompressedDataIn[1756] = 0;
decompressedDataIn[1757] = 0;
decompressedDataIn[1758] = 0;
decompressedDataIn[1759] = 0;
decompressedDataIn[1760] = 0;
decompressedDataIn[1761] = 0;
decompressedDataIn[1762] = 0;
decompressedDataIn[1763] = 0;
decompressedDataIn[1764] = 0;
decompressedDataIn[1765] = 0;
decompressedDataIn[1766] = 0;
decompressedDataIn[1767] = 0;
decompressedDataIn[1768] = 0;
decompressedDataIn[1769] = 0;
decompressedDataIn[1770] = 0;
decompressedDataIn[1771] = 0;
decompressedDataIn[1772] = 0;
decompressedDataIn[1773] = 0;
decompressedDataIn[1774] = 0;
decompressedDataIn[1775] = 0;
decompressedDataIn[1776] = 0;
decompressedDataIn[1777] = 0;
decompressedDataIn[1778] = 0;
decompressedDataIn[1779] = 0;
decompressedDataIn[1780] = 0;
decompressedDataIn[1781] = 0;
decompressedDataIn[1782] = 0;
decompressedDataIn[1783] = 0;
decompressedDataIn[1784] = 0;
decompressedDataIn[1785] = 0;
decompressedDataIn[1786] = 0;
decompressedDataIn[1787] = 0;
decompressedDataIn[1788] = 0;
decompressedDataIn[1789] = 0;
decompressedDataIn[1790] = 0;
decompressedDataIn[1791] = 0;
decompressedDataIn[1792] = 0;
decompressedDataIn[1793] = 0;
decompressedDataIn[1794] = 0;
decompressedDataIn[1795] = 0;
decompressedDataIn[1796] = 0;
decompressedDataIn[1797] = 0;
decompressedDataIn[1798] = 0;
decompressedDataIn[1799] = 0;
decompressedDataIn[1800] = 0;
decompressedDataIn[1801] = 0;
decompressedDataIn[1802] = 0;
decompressedDataIn[1803] = 0;
decompressedDataIn[1804] = 0;
decompressedDataIn[1805] = 0;
decompressedDataIn[1806] = 0;
decompressedDataIn[1807] = 0;
decompressedDataIn[1808] = 0;
decompressedDataIn[1809] = 0;
decompressedDataIn[1810] = 0;
decompressedDataIn[1811] = 0;
decompressedDataIn[1812] = 0;
decompressedDataIn[1813] = 0;
decompressedDataIn[1814] = 0;
decompressedDataIn[1815] = 0;
decompressedDataIn[1816] = 0;
decompressedDataIn[1817] = 0;
decompressedDataIn[1818] = 0;
decompressedDataIn[1819] = 0;
decompressedDataIn[1820] = 0;
decompressedDataIn[1821] = 0;
decompressedDataIn[1822] = 0;
decompressedDataIn[1823] = 0;
decompressedDataIn[1824] = 0;
decompressedDataIn[1825] = 0;
decompressedDataIn[1826] = 0;
decompressedDataIn[1827] = 0;
decompressedDataIn[1828] = 0;
decompressedDataIn[1829] = 0;
decompressedDataIn[1830] = 0;
decompressedDataIn[1831] = 0;
decompressedDataIn[1832] = 0;
decompressedDataIn[1833] = 0;
decompressedDataIn[1834] = 0;
decompressedDataIn[1835] = 0;
decompressedDataIn[1836] = 0;
decompressedDataIn[1837] = 0;
decompressedDataIn[1838] = 0;
decompressedDataIn[1839] = 0;
decompressedDataIn[1840] = 0;
decompressedDataIn[1841] = 0;
decompressedDataIn[1842] = 0;
decompressedDataIn[1843] = 0;
decompressedDataIn[1844] = 0;
decompressedDataIn[1845] = 0;
decompressedDataIn[1846] = 0;
decompressedDataIn[1847] = 0;
decompressedDataIn[1848] = 0;
decompressedDataIn[1849] = 0;
decompressedDataIn[1850] = 0;
decompressedDataIn[1851] = 0;
decompressedDataIn[1852] = 0;
decompressedDataIn[1853] = 0;
decompressedDataIn[1854] = 0;
decompressedDataIn[1855] = 0;
decompressedDataIn[1856] = 0;
decompressedDataIn[1857] = 0;
decompressedDataIn[1858] = 0;
decompressedDataIn[1859] = 0;
decompressedDataIn[1860] = 0;
decompressedDataIn[1861] = 0;
decompressedDataIn[1862] = 0;
decompressedDataIn[1863] = 0;
decompressedDataIn[1864] = 0;
decompressedDataIn[1865] = 0;
decompressedDataIn[1866] = 0;
decompressedDataIn[1867] = 0;
decompressedDataIn[1868] = 0;
decompressedDataIn[1869] = 0;
decompressedDataIn[1870] = 0;
decompressedDataIn[1871] = 0;
decompressedDataIn[1872] = 0;
decompressedDataIn[1873] = 0;
decompressedDataIn[1874] = 0;
decompressedDataIn[1875] = 0;
decompressedDataIn[1876] = 0;
decompressedDataIn[1877] = 0;
decompressedDataIn[1878] = 0;
decompressedDataIn[1879] = 0;
decompressedDataIn[1880] = 0;
decompressedDataIn[1881] = 0;
decompressedDataIn[1882] = 0;
decompressedDataIn[1883] = 0;
decompressedDataIn[1884] = 0;
decompressedDataIn[1885] = 0;
decompressedDataIn[1886] = 0;
decompressedDataIn[1887] = 0;
decompressedDataIn[1888] = 0;
decompressedDataIn[1889] = 0;
decompressedDataIn[1890] = 0;
decompressedDataIn[1891] = 0;
decompressedDataIn[1892] = 0;
decompressedDataIn[1893] = 255;
decompressedDataIn[1894] = 0;
decompressedDataIn[1895] = 0;
decompressedDataIn[1896] = 0;
decompressedDataIn[1897] = 255;
decompressedDataIn[1898] = 0;
decompressedDataIn[1899] = 0;
decompressedDataIn[1900] = 0;
decompressedDataIn[1901] = 0;
decompressedDataIn[1902] = 0;
decompressedDataIn[1903] = 255;
decompressedDataIn[1904] = 0;
decompressedDataIn[1905] = 0;
decompressedDataIn[1906] = 0;
decompressedDataIn[1907] = 0;
decompressedDataIn[1908] = 125;
decompressedDataIn[1909] = 0;
decompressedDataIn[1910] = 0;
decompressedDataIn[1911] = 0;
decompressedDataIn[1912] = 126;
decompressedDataIn[1913] = 0;
decompressedDataIn[1914] = 0;
decompressedDataIn[1915] = 0;
decompressedDataIn[1916] = 127;
decompressedDataIn[1917] = 0;
decompressedDataIn[1918] = 0;
decompressedDataIn[1919] = 0;
decompressedDataIn[1920] = 128;
decompressedDataIn[1921] = 0;
decompressedDataIn[1922] = 0;
decompressedDataIn[1923] = 0;
decompressedDataIn[1924] = 48;
decompressedDataIn[1925] = 252;
decompressedDataIn[1926] = 53;
decompressedDataIn[1927] = 247;
decompressedDataIn[1928] = 217;
decompressedDataIn[1929] = 127;
decompressedDataIn[1930] = 0;
decompressedDataIn[1931] = 0;
decompressedDataIn[1932] = 48;
decompressedDataIn[1933] = 252;
decompressedDataIn[1934] = 53;
decompressedDataIn[1935] = 247;
decompressedDataIn[1936] = 217;
decompressedDataIn[1937] = 127;
decompressedDataIn[1938] = 0;
decompressedDataIn[1939] = 0;
decompressedDataIn[1940] = 14;
decompressedDataIn[1941] = 0;
decompressedDataIn[1942] = 0;
decompressedDataIn[1943] = 0;
decompressedDataIn[1944] = 0;
decompressedDataIn[1945] = 0;
decompressedDataIn[1946] = 0;
decompressedDataIn[1947] = 0;
decompressedDataIn[1948] = 14;
decompressedDataIn[1949] = 0;
decompressedDataIn[1950] = 0;
decompressedDataIn[1951] = 0;
decompressedDataIn[1952] = 0;
decompressedDataIn[1953] = 0;
decompressedDataIn[1954] = 0;
decompressedDataIn[1955] = 0;
decompressedDataIn[1956] = 0;
decompressedDataIn[1957] = 0;
decompressedDataIn[1958] = 0;
decompressedDataIn[1959] = 0;
decompressedDataIn[1960] = 0;
decompressedDataIn[1961] = 0;
decompressedDataIn[1962] = 0;
decompressedDataIn[1963] = 0;
decompressedDataIn[1964] = 0;
decompressedDataIn[1965] = 0;
decompressedDataIn[1966] = 0;
decompressedDataIn[1967] = 0;
decompressedDataIn[1968] = 0;
decompressedDataIn[1969] = 0;
decompressedDataIn[1970] = 0;
decompressedDataIn[1971] = 0;
decompressedDataIn[1972] = 255;
decompressedDataIn[1973] = 255;
decompressedDataIn[1974] = 255;
decompressedDataIn[1975] = 255;
decompressedDataIn[1976] = 255;
decompressedDataIn[1977] = 255;
decompressedDataIn[1978] = 255;
decompressedDataIn[1979] = 255;
decompressedDataIn[1980] = 255;
decompressedDataIn[1981] = 255;
decompressedDataIn[1982] = 255;
decompressedDataIn[1983] = 255;
decompressedDataIn[1984] = 255;
decompressedDataIn[1985] = 255;
decompressedDataIn[1986] = 255;
decompressedDataIn[1987] = 255;
decompressedDataIn[1988] = 4;
decompressedDataIn[1989] = 0;
decompressedDataIn[1990] = 0;
decompressedDataIn[1991] = 0;
decompressedDataIn[1992] = 4;
decompressedDataIn[1993] = 0;
decompressedDataIn[1994] = 0;
decompressedDataIn[1995] = 0;
decompressedDataIn[1996] = 4;
decompressedDataIn[1997] = 0;
decompressedDataIn[1998] = 0;
decompressedDataIn[1999] = 0;
decompressedDataIn[2000] = 4;
decompressedDataIn[2001] = 0;
decompressedDataIn[2002] = 0;
decompressedDataIn[2003] = 0;
decompressedDataIn[2004] = 32;
decompressedDataIn[2005] = 4;
decompressedDataIn[2006] = 54;
decompressedDataIn[2007] = 247;
decompressedDataIn[2008] = 217;
decompressedDataIn[2009] = 127;
decompressedDataIn[2010] = 0;
decompressedDataIn[2011] = 0;
decompressedDataIn[2012] = 32;
decompressedDataIn[2013] = 4;
decompressedDataIn[2014] = 54;
decompressedDataIn[2015] = 247;
decompressedDataIn[2016] = 217;
decompressedDataIn[2017] = 127;
decompressedDataIn[2018] = 0;
decompressedDataIn[2019] = 0;
decompressedDataIn[2020] = 0;
decompressedDataIn[2021] = 0;
decompressedDataIn[2022] = 0;
decompressedDataIn[2023] = 0;
decompressedDataIn[2024] = 0;
decompressedDataIn[2025] = 0;
decompressedDataIn[2026] = 0;
decompressedDataIn[2027] = 0;
decompressedDataIn[2028] = 0;
decompressedDataIn[2029] = 0;
decompressedDataIn[2030] = 0;
decompressedDataIn[2031] = 0;
decompressedDataIn[2032] = 0;
decompressedDataIn[2033] = 0;
decompressedDataIn[2034] = 0;
decompressedDataIn[2035] = 0;
decompressedDataIn[2036] = 0;
decompressedDataIn[2037] = 0;
decompressedDataIn[2038] = 0;
decompressedDataIn[2039] = 0;
decompressedDataIn[2040] = 0;
decompressedDataIn[2041] = 0;
decompressedDataIn[2042] = 0;
decompressedDataIn[2043] = 0;
decompressedDataIn[2044] = 0;
decompressedDataIn[2045] = 0;
decompressedDataIn[2046] = 0;
decompressedDataIn[2047] = 0;
decompressedDataIn[2048] = 0;
decompressedDataIn[2049] = 0;
decompressedDataIn[2050] = 0;
decompressedDataIn[2051] = 0;
decompressedDataIn[2052] = 0;
decompressedDataIn[2053] = 0;
decompressedDataIn[2054] = 0;
decompressedDataIn[2055] = 0;
decompressedDataIn[2056] = 0;
decompressedDataIn[2057] = 0;
decompressedDataIn[2058] = 0;
decompressedDataIn[2059] = 0;
decompressedDataIn[2060] = 0;
decompressedDataIn[2061] = 0;
decompressedDataIn[2062] = 0;
decompressedDataIn[2063] = 0;
decompressedDataIn[2064] = 0;
decompressedDataIn[2065] = 0;
decompressedDataIn[2066] = 0;
decompressedDataIn[2067] = 0;
decompressedDataIn[2068] = 0;
decompressedDataIn[2069] = 0;
decompressedDataIn[2070] = 0;
decompressedDataIn[2071] = 0;
decompressedDataIn[2072] = 0;
decompressedDataIn[2073] = 0;
decompressedDataIn[2074] = 0;
decompressedDataIn[2075] = 0;
decompressedDataIn[2076] = 0;
decompressedDataIn[2077] = 0;
decompressedDataIn[2078] = 0;
decompressedDataIn[2079] = 0;
decompressedDataIn[2080] = 0;
decompressedDataIn[2081] = 0;
decompressedDataIn[2082] = 0;
decompressedDataIn[2083] = 0;
decompressedDataIn[2084] = 0;
decompressedDataIn[2085] = 0;
decompressedDataIn[2086] = 0;
decompressedDataIn[2087] = 0;
decompressedDataIn[2088] = 0;
decompressedDataIn[2089] = 0;
decompressedDataIn[2090] = 0;
decompressedDataIn[2091] = 0;
decompressedDataIn[2092] = 0;
decompressedDataIn[2093] = 0;
decompressedDataIn[2094] = 0;
decompressedDataIn[2095] = 0;
decompressedDataIn[2096] = 0;
decompressedDataIn[2097] = 0;
decompressedDataIn[2098] = 0;
decompressedDataIn[2099] = 0;
decompressedDataIn[2100] = 0;
decompressedDataIn[2101] = 0;
decompressedDataIn[2102] = 0;
decompressedDataIn[2103] = 0;
decompressedDataIn[2104] = 0;
decompressedDataIn[2105] = 0;
decompressedDataIn[2106] = 0;
decompressedDataIn[2107] = 0;
decompressedDataIn[2108] = 0;
decompressedDataIn[2109] = 0;
decompressedDataIn[2110] = 0;
decompressedDataIn[2111] = 0;
decompressedDataIn[2112] = 0;
decompressedDataIn[2113] = 0;
decompressedDataIn[2114] = 0;
decompressedDataIn[2115] = 0;
decompressedDataIn[2116] = 0;
decompressedDataIn[2117] = 0;
decompressedDataIn[2118] = 0;
decompressedDataIn[2119] = 0;
decompressedDataIn[2120] = 0;
decompressedDataIn[2121] = 0;
decompressedDataIn[2122] = 0;
decompressedDataIn[2123] = 0;
decompressedDataIn[2124] = 0;
decompressedDataIn[2125] = 0;
decompressedDataIn[2126] = 0;
decompressedDataIn[2127] = 0;
decompressedDataIn[2128] = 0;
decompressedDataIn[2129] = 0;
decompressedDataIn[2130] = 0;
decompressedDataIn[2131] = 0;
decompressedDataIn[2132] = 155;
decompressedDataIn[2133] = 80;
decompressedDataIn[2134] = 214;
decompressedDataIn[2135] = 97;
decompressedDataIn[2136] = 58;
decompressedDataIn[2137] = 127;
decompressedDataIn[2138] = 0;
decompressedDataIn[2139] = 0;
decompressedDataIn[2140] = 10;
decompressedDataIn[2141] = 0;
decompressedDataIn[2142] = 0;
decompressedDataIn[2143] = 0;
decompressedDataIn[2144] = 0;
decompressedDataIn[2145] = 0;
decompressedDataIn[2146] = 0;
decompressedDataIn[2147] = 0;
decompressedDataIn[2148] = 0;
decompressedDataIn[2149] = 0;
decompressedDataIn[2150] = 0;
decompressedDataIn[2151] = 0;
decompressedDataIn[2152] = 0;
decompressedDataIn[2153] = 85;
decompressedDataIn[2154] = 0;
decompressedDataIn[2155] = 0;
decompressedDataIn[2156] = 0;
decompressedDataIn[2157] = 0;
decompressedDataIn[2158] = 0;
decompressedDataIn[2159] = 0;
decompressedDataIn[2160] = 0;
decompressedDataIn[2161] = 0;
decompressedDataIn[2162] = 0;
decompressedDataIn[2163] = 0;
decompressedDataIn[2164] = 170;
decompressedDataIn[2165] = 80;
decompressedDataIn[2166] = 214;
decompressedDataIn[2167] = 97;
decompressedDataIn[2168] = 58;
decompressedDataIn[2169] = 127;
decompressedDataIn[2170] = 0;
decompressedDataIn[2171] = 0;
decompressedDataIn[2172] = 11;
decompressedDataIn[2173] = 0;
decompressedDataIn[2174] = 0;
decompressedDataIn[2175] = 0;
decompressedDataIn[2176] = 0;
decompressedDataIn[2177] = 0;
decompressedDataIn[2178] = 0;
decompressedDataIn[2179] = 0;
decompressedDataIn[2180] = 0;
decompressedDataIn[2181] = 0;
decompressedDataIn[2182] = 0;
decompressedDataIn[2183] = 0;
decompressedDataIn[2184] = 0;
decompressedDataIn[2185] = 85;
decompressedDataIn[2186] = 0;
decompressedDataIn[2187] = 0;
decompressedDataIn[2188] = 0;
decompressedDataIn[2189] = 0;
decompressedDataIn[2190] = 0;
decompressedDataIn[2191] = 0;
decompressedDataIn[2192] = 0;
decompressedDataIn[2193] = 0;
decompressedDataIn[2194] = 0;
decompressedDataIn[2195] = 0;
decompressedDataIn[2196] = 180;
decompressedDataIn[2197] = 80;
decompressedDataIn[2198] = 214;
decompressedDataIn[2199] = 97;
decompressedDataIn[2200] = 58;
decompressedDataIn[2201] = 127;
decompressedDataIn[2202] = 0;
decompressedDataIn[2203] = 0;
decompressedDataIn[2204] = 8;
decompressedDataIn[2205] = 0;
decompressedDataIn[2206] = 0;
decompressedDataIn[2207] = 0;
decompressedDataIn[2208] = 0;
decompressedDataIn[2209] = 0;
decompressedDataIn[2210] = 0;
decompressedDataIn[2211] = 0;
decompressedDataIn[2212] = 0;
decompressedDataIn[2213] = 0;
decompressedDataIn[2214] = 0;
decompressedDataIn[2215] = 0;
decompressedDataIn[2216] = 0;
decompressedDataIn[2217] = 85;
decompressedDataIn[2218] = 0;
decompressedDataIn[2219] = 0;
decompressedDataIn[2220] = 0;
decompressedDataIn[2221] = 0;
decompressedDataIn[2222] = 0;
decompressedDataIn[2223] = 0;
decompressedDataIn[2224] = 0;
decompressedDataIn[2225] = 0;
decompressedDataIn[2226] = 0;
decompressedDataIn[2227] = 0;
decompressedDataIn[2228] = 6;
decompressedDataIn[2229] = 0;
decompressedDataIn[2230] = 0;
decompressedDataIn[2231] = 0;
decompressedDataIn[2232] = 64;
decompressedDataIn[2233] = 4;
decompressedDataIn[2234] = 0;
decompressedDataIn[2235] = 0;
decompressedDataIn[2236] = 2;
decompressedDataIn[2237] = 2;
decompressedDataIn[2238] = 0;
decompressedDataIn[2239] = 0;
decompressedDataIn[2240] = 76;
decompressedDataIn[2241] = 73;
decompressedDataIn[2242] = 78;
decompressedDataIn[2243] = 85;
decompressedDataIn[2244] = 88;
decompressedDataIn[2245] = 0;
decompressedDataIn[2246] = 0;
decompressedDataIn[2247] = 0;
decompressedDataIn[2248] = 255;
decompressedDataIn[2249] = 255;
decompressedDataIn[2250] = 255;
decompressedDataIn[2251] = 255;
decompressedDataIn[2252] = 255;
decompressedDataIn[2253] = 0;
decompressedDataIn[2254] = 255;
decompressedDataIn[2255] = 7;
decompressedDataIn[2256] = 106;
decompressedDataIn[2257] = 102;
decompressedDataIn[2258] = 14;
decompressedDataIn[2259] = 210;
decompressedDataIn[2260] = 225;
decompressedDataIn[2261] = 85;
decompressedDataIn[2262] = 0;
decompressedDataIn[2263] = 0;
decompressedDataIn[2264] = 0;
decompressedDataIn[2265] = 194;
decompressedDataIn[2266] = 55;
decompressedDataIn[2267] = 75;
decompressedDataIn[2268] = 254;
decompressedDataIn[2269] = 127;
decompressedDataIn[2270] = 0;
decompressedDataIn[2271] = 0;
decompressedDataIn[2272] = 160;
decompressedDataIn[2273] = 31;
decompressedDataIn[2274] = 0;
decompressedDataIn[2275] = 0;
    $display("testing");
decompressedDataIn[2276] = 0;
decompressedDataIn[2277] = 0;
decompressedDataIn[2278] = 0;
decompressedDataIn[2279] = 0;
decompressedDataIn[2280] = 0;
decompressedDataIn[2281] = 0;
decompressedDataIn[2282] = 0;
decompressedDataIn[2283] = 0;
decompressedDataIn[2284] = 0;
decompressedDataIn[2285] = 0;
decompressedDataIn[2286] = 0;
decompressedDataIn[2287] = 0;
decompressedDataIn[2288] = 0;
decompressedDataIn[2289] = 0;
decompressedDataIn[2290] = 0;
decompressedDataIn[2291] = 0;
decompressedDataIn[2292] = 0;
decompressedDataIn[2293] = 0;
decompressedDataIn[2294] = 0;
decompressedDataIn[2295] = 0;
decompressedDataIn[2296] = 0;
decompressedDataIn[2297] = 0;
decompressedDataIn[2298] = 0;
decompressedDataIn[2299] = 0;
decompressedDataIn[2300] = 0;
decompressedDataIn[2301] = 0;
decompressedDataIn[2302] = 0;
decompressedDataIn[2303] = 0;
decompressedDataIn[2304] = 0;
decompressedDataIn[2305] = 0;
decompressedDataIn[2306] = 0;
decompressedDataIn[2307] = 0;
decompressedDataIn[2308] = 0;
decompressedDataIn[2309] = 0;
decompressedDataIn[2310] = 0;
decompressedDataIn[2311] = 0;
decompressedDataIn[2312] = 0;
decompressedDataIn[2313] = 0;
decompressedDataIn[2314] = 0;
decompressedDataIn[2315] = 0;
decompressedDataIn[2316] = 0;
decompressedDataIn[2317] = 0;
decompressedDataIn[2318] = 0;
decompressedDataIn[2319] = 0;
decompressedDataIn[2320] = 0;
decompressedDataIn[2321] = 0;
decompressedDataIn[2322] = 0;
decompressedDataIn[2323] = 0;
decompressedDataIn[2324] = 0;
decompressedDataIn[2325] = 0;
decompressedDataIn[2326] = 0;
decompressedDataIn[2327] = 0;
decompressedDataIn[2328] = 0;
decompressedDataIn[2329] = 0;
decompressedDataIn[2330] = 0;
decompressedDataIn[2331] = 0;
decompressedDataIn[2332] = 0;
decompressedDataIn[2333] = 0;
decompressedDataIn[2334] = 0;
decompressedDataIn[2335] = 0;
decompressedDataIn[2336] = 0;
decompressedDataIn[2337] = 0;
decompressedDataIn[2338] = 0;
decompressedDataIn[2339] = 0;
decompressedDataIn[2340] = 0;
decompressedDataIn[2341] = 0;
decompressedDataIn[2342] = 0;
decompressedDataIn[2343] = 0;
decompressedDataIn[2344] = 0;
decompressedDataIn[2345] = 0;
decompressedDataIn[2346] = 0;
decompressedDataIn[2347] = 0;
decompressedDataIn[2348] = 0;
decompressedDataIn[2349] = 0;
decompressedDataIn[2350] = 0;
decompressedDataIn[2351] = 0;
decompressedDataIn[2352] = 0;
decompressedDataIn[2353] = 0;
decompressedDataIn[2354] = 0;
decompressedDataIn[2355] = 0;
decompressedDataIn[2356] = 0;
decompressedDataIn[2357] = 0;
decompressedDataIn[2358] = 0;
decompressedDataIn[2359] = 0;
decompressedDataIn[2360] = 0;
decompressedDataIn[2361] = 0;
decompressedDataIn[2362] = 0;
decompressedDataIn[2363] = 0;
decompressedDataIn[2364] = 0;
decompressedDataIn[2365] = 0;
decompressedDataIn[2366] = 0;
decompressedDataIn[2367] = 0;
decompressedDataIn[2368] = 0;
decompressedDataIn[2369] = 0;
decompressedDataIn[2370] = 0;
decompressedDataIn[2371] = 0;
decompressedDataIn[2372] = 0;
decompressedDataIn[2373] = 0;
decompressedDataIn[2374] = 0;
decompressedDataIn[2375] = 0;
decompressedDataIn[2376] = 0;
decompressedDataIn[2377] = 0;
decompressedDataIn[2378] = 0;
decompressedDataIn[2379] = 0;
decompressedDataIn[2380] = 0;
decompressedDataIn[2381] = 0;
decompressedDataIn[2382] = 0;
decompressedDataIn[2383] = 0;
decompressedDataIn[2384] = 0;
decompressedDataIn[2385] = 0;
decompressedDataIn[2386] = 0;
decompressedDataIn[2387] = 0;
decompressedDataIn[2388] = 0;
decompressedDataIn[2389] = 0;
decompressedDataIn[2390] = 0;
decompressedDataIn[2391] = 0;
decompressedDataIn[2392] = 0;
decompressedDataIn[2393] = 0;
decompressedDataIn[2394] = 0;
decompressedDataIn[2395] = 0;
decompressedDataIn[2396] = 0;
decompressedDataIn[2397] = 0;
decompressedDataIn[2398] = 0;
decompressedDataIn[2399] = 0;
decompressedDataIn[2400] = 0;
decompressedDataIn[2401] = 0;
decompressedDataIn[2402] = 0;
decompressedDataIn[2403] = 0;
decompressedDataIn[2404] = 0;
decompressedDataIn[2405] = 0;
decompressedDataIn[2406] = 0;
decompressedDataIn[2407] = 0;
decompressedDataIn[2408] = 0;
decompressedDataIn[2409] = 0;
decompressedDataIn[2410] = 0;
decompressedDataIn[2411] = 0;
decompressedDataIn[2412] = 0;
decompressedDataIn[2413] = 0;
decompressedDataIn[2414] = 0;
decompressedDataIn[2415] = 0;
decompressedDataIn[2416] = 0;
decompressedDataIn[2417] = 0;
decompressedDataIn[2418] = 0;
decompressedDataIn[2419] = 0;
decompressedDataIn[2420] = 0;
decompressedDataIn[2421] = 0;
decompressedDataIn[2422] = 0;
decompressedDataIn[2423] = 0;
decompressedDataIn[2424] = 0;
decompressedDataIn[2425] = 255;
decompressedDataIn[2426] = 0;
decompressedDataIn[2427] = 0;
decompressedDataIn[2428] = 0;
decompressedDataIn[2429] = 255;
decompressedDataIn[2430] = 0;
decompressedDataIn[2431] = 0;
decompressedDataIn[2432] = 0;
decompressedDataIn[2433] = 0;
decompressedDataIn[2434] = 0;
decompressedDataIn[2435] = 255;
decompressedDataIn[2436] = 0;
decompressedDataIn[2437] = 0;
decompressedDataIn[2438] = 0;
decompressedDataIn[2439] = 0;
decompressedDataIn[2440] = 125;
decompressedDataIn[2441] = 0;
decompressedDataIn[2442] = 0;
decompressedDataIn[2443] = 0;
decompressedDataIn[2444] = 126;
decompressedDataIn[2445] = 0;
decompressedDataIn[2446] = 0;
decompressedDataIn[2447] = 0;
decompressedDataIn[2448] = 127;
decompressedDataIn[2449] = 0;
decompressedDataIn[2450] = 0;
decompressedDataIn[2451] = 0;
decompressedDataIn[2452] = 128;
decompressedDataIn[2453] = 0;
decompressedDataIn[2454] = 0;
decompressedDataIn[2455] = 0;
decompressedDataIn[2456] = 48;
decompressedDataIn[2457] = 252;
decompressedDataIn[2458] = 53;
decompressedDataIn[2459] = 247;
decompressedDataIn[2460] = 217;
decompressedDataIn[2461] = 127;
decompressedDataIn[2462] = 0;
decompressedDataIn[2463] = 0;
decompressedDataIn[2464] = 48;
decompressedDataIn[2465] = 252;
decompressedDataIn[2466] = 53;
decompressedDataIn[2467] = 247;
decompressedDataIn[2468] = 217;
decompressedDataIn[2469] = 127;
decompressedDataIn[2470] = 0;
decompressedDataIn[2471] = 0;
decompressedDataIn[2472] = 14;
decompressedDataIn[2473] = 0;
decompressedDataIn[2474] = 0;
decompressedDataIn[2475] = 0;
decompressedDataIn[2476] = 0;
decompressedDataIn[2477] = 0;
decompressedDataIn[2478] = 0;
decompressedDataIn[2479] = 0;
decompressedDataIn[2480] = 14;
decompressedDataIn[2481] = 0;
decompressedDataIn[2482] = 0;
decompressedDataIn[2483] = 0;
decompressedDataIn[2484] = 0;
decompressedDataIn[2485] = 0;
decompressedDataIn[2486] = 0;
decompressedDataIn[2487] = 0;
decompressedDataIn[2488] = 0;
decompressedDataIn[2489] = 0;
decompressedDataIn[2490] = 0;
decompressedDataIn[2491] = 0;
decompressedDataIn[2492] = 0;
decompressedDataIn[2493] = 0;
decompressedDataIn[2494] = 0;
decompressedDataIn[2495] = 0;
decompressedDataIn[2496] = 0;
decompressedDataIn[2497] = 0;
decompressedDataIn[2498] = 0;
decompressedDataIn[2499] = 0;
decompressedDataIn[2500] = 0;
decompressedDataIn[2501] = 0;
decompressedDataIn[2502] = 0;
decompressedDataIn[2503] = 0;
decompressedDataIn[2504] = 255;
decompressedDataIn[2505] = 255;
decompressedDataIn[2506] = 255;
decompressedDataIn[2507] = 255;
decompressedDataIn[2508] = 255;
decompressedDataIn[2509] = 255;
decompressedDataIn[2510] = 255;
decompressedDataIn[2511] = 255;
decompressedDataIn[2512] = 255;
decompressedDataIn[2513] = 255;
decompressedDataIn[2514] = 255;
decompressedDataIn[2515] = 255;
decompressedDataIn[2516] = 255;
decompressedDataIn[2517] = 255;
decompressedDataIn[2518] = 255;
decompressedDataIn[2519] = 255;
decompressedDataIn[2520] = 4;
decompressedDataIn[2521] = 0;
decompressedDataIn[2522] = 0;
decompressedDataIn[2523] = 0;
decompressedDataIn[2524] = 4;
decompressedDataIn[2525] = 0;
decompressedDataIn[2526] = 0;
decompressedDataIn[2527] = 0;
decompressedDataIn[2528] = 4;
decompressedDataIn[2529] = 0;
decompressedDataIn[2530] = 0;
decompressedDataIn[2531] = 0;
decompressedDataIn[2532] = 4;
decompressedDataIn[2533] = 0;
decompressedDataIn[2534] = 0;
decompressedDataIn[2535] = 0;
decompressedDataIn[2536] = 32;
decompressedDataIn[2537] = 4;
decompressedDataIn[2538] = 54;
decompressedDataIn[2539] = 247;
decompressedDataIn[2540] = 217;
decompressedDataIn[2541] = 127;
decompressedDataIn[2542] = 0;
decompressedDataIn[2543] = 0;
decompressedDataIn[2544] = 32;
decompressedDataIn[2545] = 4;
decompressedDataIn[2546] = 54;
decompressedDataIn[2547] = 247;
decompressedDataIn[2548] = 217;
decompressedDataIn[2549] = 127;
decompressedDataIn[2550] = 0;
decompressedDataIn[2551] = 0;
decompressedDataIn[2552] = 0;
decompressedDataIn[2553] = 0;
decompressedDataIn[2554] = 0;
decompressedDataIn[2555] = 0;
decompressedDataIn[2556] = 0;
decompressedDataIn[2557] = 0;
decompressedDataIn[2558] = 0;
decompressedDataIn[2559] = 0;
decompressedDataIn[2560] = 0;
decompressedDataIn[2561] = 0;
decompressedDataIn[2562] = 0;
decompressedDataIn[2563] = 0;
decompressedDataIn[2564] = 0;
decompressedDataIn[2565] = 0;
decompressedDataIn[2566] = 0;
decompressedDataIn[2567] = 0;
decompressedDataIn[2568] = 0;
decompressedDataIn[2569] = 0;
decompressedDataIn[2570] = 0;
decompressedDataIn[2571] = 0;
decompressedDataIn[2572] = 0;
decompressedDataIn[2573] = 0;
decompressedDataIn[2574] = 0;
decompressedDataIn[2575] = 0;
decompressedDataIn[2576] = 0;
decompressedDataIn[2577] = 0;
decompressedDataIn[2578] = 0;
decompressedDataIn[2579] = 0;
decompressedDataIn[2580] = 0;
decompressedDataIn[2581] = 0;
decompressedDataIn[2582] = 0;
decompressedDataIn[2583] = 0;
decompressedDataIn[2584] = 0;
decompressedDataIn[2585] = 0;
decompressedDataIn[2586] = 0;
decompressedDataIn[2587] = 0;
decompressedDataIn[2588] = 0;
decompressedDataIn[2589] = 0;
decompressedDataIn[2590] = 0;
decompressedDataIn[2591] = 0;
decompressedDataIn[2592] = 0;
decompressedDataIn[2593] = 0;
decompressedDataIn[2594] = 0;
decompressedDataIn[2595] = 0;
decompressedDataIn[2596] = 0;
decompressedDataIn[2597] = 0;
decompressedDataIn[2598] = 0;
decompressedDataIn[2599] = 0;
decompressedDataIn[2600] = 0;
decompressedDataIn[2601] = 0;
decompressedDataIn[2602] = 0;
decompressedDataIn[2603] = 0;
decompressedDataIn[2604] = 0;
decompressedDataIn[2605] = 0;
decompressedDataIn[2606] = 0;
decompressedDataIn[2607] = 0;
decompressedDataIn[2608] = 0;
decompressedDataIn[2609] = 0;
decompressedDataIn[2610] = 0;
decompressedDataIn[2611] = 0;
decompressedDataIn[2612] = 0;
decompressedDataIn[2613] = 0;
decompressedDataIn[2614] = 0;
decompressedDataIn[2615] = 0;
decompressedDataIn[2616] = 0;
decompressedDataIn[2617] = 0;
decompressedDataIn[2618] = 0;
decompressedDataIn[2619] = 0;
decompressedDataIn[2620] = 0;
decompressedDataIn[2621] = 0;
decompressedDataIn[2622] = 0;
decompressedDataIn[2623] = 0;
decompressedDataIn[2624] = 0;
decompressedDataIn[2625] = 0;
decompressedDataIn[2626] = 0;
decompressedDataIn[2627] = 0;
decompressedDataIn[2628] = 0;
decompressedDataIn[2629] = 0;
decompressedDataIn[2630] = 0;
decompressedDataIn[2631] = 0;
decompressedDataIn[2632] = 0;
decompressedDataIn[2633] = 0;
decompressedDataIn[2634] = 0;
decompressedDataIn[2635] = 0;
decompressedDataIn[2636] = 0;
decompressedDataIn[2637] = 0;
decompressedDataIn[2638] = 0;
decompressedDataIn[2639] = 0;
decompressedDataIn[2640] = 0;
decompressedDataIn[2641] = 0;
decompressedDataIn[2642] = 0;
decompressedDataIn[2643] = 0;
decompressedDataIn[2644] = 0;
decompressedDataIn[2645] = 0;
decompressedDataIn[2646] = 0;
decompressedDataIn[2647] = 0;
decompressedDataIn[2648] = 0;
decompressedDataIn[2649] = 0;
decompressedDataIn[2650] = 0;
decompressedDataIn[2651] = 0;
decompressedDataIn[2652] = 0;
decompressedDataIn[2653] = 0;
decompressedDataIn[2654] = 0;
decompressedDataIn[2655] = 0;
decompressedDataIn[2656] = 0;
decompressedDataIn[2657] = 0;
decompressedDataIn[2658] = 0;
decompressedDataIn[2659] = 0;
decompressedDataIn[2660] = 0;
decompressedDataIn[2661] = 0;
decompressedDataIn[2662] = 0;
decompressedDataIn[2663] = 0;
decompressedDataIn[2664] = 0;
decompressedDataIn[2665] = 0;
decompressedDataIn[2666] = 0;
decompressedDataIn[2667] = 0;
decompressedDataIn[2668] = 0;
decompressedDataIn[2669] = 0;
decompressedDataIn[2670] = 0;
decompressedDataIn[2671] = 0;
decompressedDataIn[2672] = 0;
decompressedDataIn[2673] = 0;
decompressedDataIn[2674] = 0;
decompressedDataIn[2675] = 0;
decompressedDataIn[2676] = 0;
decompressedDataIn[2677] = 0;
decompressedDataIn[2678] = 0;
decompressedDataIn[2679] = 0;
decompressedDataIn[2680] = 0;
decompressedDataIn[2681] = 0;
decompressedDataIn[2682] = 0;
decompressedDataIn[2683] = 0;
decompressedDataIn[2684] = 0;
decompressedDataIn[2685] = 0;
decompressedDataIn[2686] = 0;
decompressedDataIn[2687] = 0;
decompressedDataIn[2688] = 0;
decompressedDataIn[2689] = 0;
decompressedDataIn[2690] = 0;
decompressedDataIn[2691] = 0;
decompressedDataIn[2692] = 0;
decompressedDataIn[2693] = 0;
decompressedDataIn[2694] = 0;
decompressedDataIn[2695] = 0;
decompressedDataIn[2696] = 0;
decompressedDataIn[2697] = 0;
decompressedDataIn[2698] = 0;
decompressedDataIn[2699] = 0;
decompressedDataIn[2700] = 0;
decompressedDataIn[2701] = 0;
decompressedDataIn[2702] = 0;
decompressedDataIn[2703] = 0;
decompressedDataIn[2704] = 0;
decompressedDataIn[2705] = 0;
decompressedDataIn[2706] = 0;
decompressedDataIn[2707] = 0;
decompressedDataIn[2708] = 0;
decompressedDataIn[2709] = 0;
decompressedDataIn[2710] = 0;
decompressedDataIn[2711] = 0;
decompressedDataIn[2712] = 31;
decompressedDataIn[2713] = 0;
decompressedDataIn[2714] = 0;
decompressedDataIn[2715] = 0;
decompressedDataIn[2716] = 0;
decompressedDataIn[2717] = 0;
decompressedDataIn[2718] = 0;
decompressedDataIn[2719] = 0;
decompressedDataIn[2720] = 0;
decompressedDataIn[2721] = 0;
decompressedDataIn[2722] = 0;
decompressedDataIn[2723] = 0;
decompressedDataIn[2724] = 0;
decompressedDataIn[2725] = 0;
decompressedDataIn[2726] = 0;
decompressedDataIn[2727] = 0;
decompressedDataIn[2728] = 0;
decompressedDataIn[2729] = 0;
decompressedDataIn[2730] = 0;
decompressedDataIn[2731] = 0;
decompressedDataIn[2732] = 0;
decompressedDataIn[2733] = 0;
decompressedDataIn[2734] = 0;
decompressedDataIn[2735] = 0;
decompressedDataIn[2736] = 0;
decompressedDataIn[2737] = 0;
decompressedDataIn[2738] = 0;
decompressedDataIn[2739] = 0;
decompressedDataIn[2740] = 0;
decompressedDataIn[2741] = 0;
decompressedDataIn[2742] = 0;
decompressedDataIn[2743] = 0;
decompressedDataIn[2744] = 0;
decompressedDataIn[2745] = 0;
decompressedDataIn[2746] = 0;
decompressedDataIn[2747] = 0;
decompressedDataIn[2748] = 0;
decompressedDataIn[2749] = 0;
decompressedDataIn[2750] = 0;
decompressedDataIn[2751] = 0;
decompressedDataIn[2752] = 0;
decompressedDataIn[2753] = 0;
decompressedDataIn[2754] = 0;
decompressedDataIn[2755] = 0;
decompressedDataIn[2756] = 0;
decompressedDataIn[2757] = 0;
decompressedDataIn[2758] = 0;
decompressedDataIn[2759] = 0;
decompressedDataIn[2760] = 31;
decompressedDataIn[2761] = 0;
decompressedDataIn[2762] = 0;
decompressedDataIn[2763] = 0;
decompressedDataIn[2764] = 0;
decompressedDataIn[2765] = 0;
decompressedDataIn[2766] = 0;
decompressedDataIn[2767] = 0;
decompressedDataIn[2768] = 0;
decompressedDataIn[2769] = 0;
decompressedDataIn[2770] = 0;
decompressedDataIn[2771] = 0;
decompressedDataIn[2772] = 0;
decompressedDataIn[2773] = 0;
decompressedDataIn[2774] = 0;
decompressedDataIn[2775] = 0;
decompressedDataIn[2776] = 0;
decompressedDataIn[2777] = 0;
decompressedDataIn[2778] = 0;
decompressedDataIn[2779] = 0;
decompressedDataIn[2780] = 0;
decompressedDataIn[2781] = 0;
decompressedDataIn[2782] = 0;
decompressedDataIn[2783] = 0;
decompressedDataIn[2784] = 0;
decompressedDataIn[2785] = 0;
decompressedDataIn[2786] = 0;
decompressedDataIn[2787] = 0;
decompressedDataIn[2788] = 0;
decompressedDataIn[2789] = 0;
decompressedDataIn[2790] = 0;
decompressedDataIn[2791] = 0;
decompressedDataIn[2792] = 0;
decompressedDataIn[2793] = 0;
decompressedDataIn[2794] = 0;
decompressedDataIn[2795] = 0;
decompressedDataIn[2796] = 0;
decompressedDataIn[2797] = 0;
decompressedDataIn[2798] = 0;
decompressedDataIn[2799] = 0;
decompressedDataIn[2800] = 0;
decompressedDataIn[2801] = 0;
decompressedDataIn[2802] = 0;
decompressedDataIn[2803] = 0;
decompressedDataIn[2804] = 0;
decompressedDataIn[2805] = 0;
decompressedDataIn[2806] = 0;
decompressedDataIn[2807] = 0;
decompressedDataIn[2808] = 0;
decompressedDataIn[2809] = 0;
decompressedDataIn[2810] = 0;
decompressedDataIn[2811] = 0;
decompressedDataIn[2812] = 0;
decompressedDataIn[2813] = 0;
decompressedDataIn[2814] = 0;
decompressedDataIn[2815] = 0;
decompressedDataIn[2816] = 0;
decompressedDataIn[2817] = 0;
decompressedDataIn[2818] = 0;
decompressedDataIn[2819] = 0;
decompressedDataIn[2820] = 0;
decompressedDataIn[2821] = 0;
decompressedDataIn[2822] = 0;
decompressedDataIn[2823] = 0;
decompressedDataIn[2824] = 0;
decompressedDataIn[2825] = 0;
decompressedDataIn[2826] = 0;
decompressedDataIn[2827] = 0;
decompressedDataIn[2828] = 0;
decompressedDataIn[2829] = 0;
decompressedDataIn[2830] = 0;
decompressedDataIn[2831] = 0;
decompressedDataIn[2832] = 0;
decompressedDataIn[2833] = 0;
decompressedDataIn[2834] = 0;
decompressedDataIn[2835] = 0;
decompressedDataIn[2836] = 0;
decompressedDataIn[2837] = 0;
decompressedDataIn[2838] = 0;
decompressedDataIn[2839] = 0;
decompressedDataIn[2840] = 0;
decompressedDataIn[2841] = 0;
decompressedDataIn[2842] = 0;
decompressedDataIn[2843] = 0;
decompressedDataIn[2844] = 0;
decompressedDataIn[2845] = 0;
decompressedDataIn[2846] = 0;
decompressedDataIn[2847] = 0;
decompressedDataIn[2848] = 0;
decompressedDataIn[2849] = 0;
decompressedDataIn[2850] = 0;
decompressedDataIn[2851] = 0;
decompressedDataIn[2852] = 0;
decompressedDataIn[2853] = 0;
decompressedDataIn[2854] = 0;
decompressedDataIn[2855] = 0;
decompressedDataIn[2856] = 0;
decompressedDataIn[2857] = 0;
decompressedDataIn[2858] = 0;
decompressedDataIn[2859] = 0;
decompressedDataIn[2860] = 0;
decompressedDataIn[2861] = 0;
decompressedDataIn[2862] = 0;
decompressedDataIn[2863] = 0;
decompressedDataIn[2864] = 0;
decompressedDataIn[2865] = 0;
decompressedDataIn[2866] = 0;
decompressedDataIn[2867] = 0;
decompressedDataIn[2868] = 0;
decompressedDataIn[2869] = 0;
decompressedDataIn[2870] = 0;
decompressedDataIn[2871] = 0;
decompressedDataIn[2872] = 0;
decompressedDataIn[2873] = 0;
decompressedDataIn[2874] = 0;
decompressedDataIn[2875] = 0;
decompressedDataIn[2876] = 0;
decompressedDataIn[2877] = 0;
decompressedDataIn[2878] = 0;
decompressedDataIn[2879] = 0;
decompressedDataIn[2880] = 0;
decompressedDataIn[2881] = 0;
decompressedDataIn[2882] = 0;
decompressedDataIn[2883] = 0;
decompressedDataIn[2884] = 0;
decompressedDataIn[2885] = 0;
decompressedDataIn[2886] = 0;
decompressedDataIn[2887] = 0;
decompressedDataIn[2888] = 0;
decompressedDataIn[2889] = 0;
decompressedDataIn[2890] = 0;
decompressedDataIn[2891] = 0;
decompressedDataIn[2892] = 0;
decompressedDataIn[2893] = 0;
decompressedDataIn[2894] = 0;
decompressedDataIn[2895] = 0;
decompressedDataIn[2896] = 0;
decompressedDataIn[2897] = 0;
decompressedDataIn[2898] = 0;
decompressedDataIn[2899] = 0;
decompressedDataIn[2900] = 0;
decompressedDataIn[2901] = 0;
decompressedDataIn[2902] = 0;
decompressedDataIn[2903] = 0;
decompressedDataIn[2904] = 0;
decompressedDataIn[2905] = 0;
decompressedDataIn[2906] = 0;
decompressedDataIn[2907] = 0;
decompressedDataIn[2908] = 0;
decompressedDataIn[2909] = 0;
decompressedDataIn[2910] = 0;
decompressedDataIn[2911] = 0;
decompressedDataIn[2912] = 0;
decompressedDataIn[2913] = 0;
decompressedDataIn[2914] = 0;
decompressedDataIn[2915] = 0;
decompressedDataIn[2916] = 0;
decompressedDataIn[2917] = 0;
decompressedDataIn[2918] = 0;
decompressedDataIn[2919] = 0;
decompressedDataIn[2920] = 0;
decompressedDataIn[2921] = 0;
decompressedDataIn[2922] = 0;
decompressedDataIn[2923] = 0;
decompressedDataIn[2924] = 0;
decompressedDataIn[2925] = 0;
decompressedDataIn[2926] = 0;
decompressedDataIn[2927] = 0;
decompressedDataIn[2928] = 0;
decompressedDataIn[2929] = 0;
decompressedDataIn[2930] = 0;
decompressedDataIn[2931] = 0;
decompressedDataIn[2932] = 0;
decompressedDataIn[2933] = 0;
decompressedDataIn[2934] = 0;
decompressedDataIn[2935] = 0;
decompressedDataIn[2936] = 0;
decompressedDataIn[2937] = 0;
decompressedDataIn[2938] = 0;
decompressedDataIn[2939] = 0;
decompressedDataIn[2940] = 0;
decompressedDataIn[2941] = 0;
decompressedDataIn[2942] = 0;
decompressedDataIn[2943] = 0;
decompressedDataIn[2944] = 0;
decompressedDataIn[2945] = 0;
decompressedDataIn[2946] = 0;
decompressedDataIn[2947] = 0;
decompressedDataIn[2948] = 0;
decompressedDataIn[2949] = 0;
decompressedDataIn[2950] = 0;
decompressedDataIn[2951] = 0;
decompressedDataIn[2952] = 0;
decompressedDataIn[2953] = 0;
decompressedDataIn[2954] = 0;
decompressedDataIn[2955] = 0;
decompressedDataIn[2956] = 0;
decompressedDataIn[2957] = 0;
decompressedDataIn[2958] = 0;
decompressedDataIn[2959] = 0;
decompressedDataIn[2960] = 0;
decompressedDataIn[2961] = 0;
decompressedDataIn[2962] = 0;
decompressedDataIn[2963] = 0;
decompressedDataIn[2964] = 0;
decompressedDataIn[2965] = 0;
decompressedDataIn[2966] = 0;
decompressedDataIn[2967] = 0;
decompressedDataIn[2968] = 0;
decompressedDataIn[2969] = 0;
decompressedDataIn[2970] = 0;
decompressedDataIn[2971] = 0;
decompressedDataIn[2972] = 0;
decompressedDataIn[2973] = 0;
decompressedDataIn[2974] = 0;
decompressedDataIn[2975] = 0;
decompressedDataIn[2976] = 0;
decompressedDataIn[2977] = 0;
decompressedDataIn[2978] = 0;
decompressedDataIn[2979] = 0;
decompressedDataIn[2980] = 0;
decompressedDataIn[2981] = 0;
decompressedDataIn[2982] = 0;
decompressedDataIn[2983] = 0;
decompressedDataIn[2984] = 0;
decompressedDataIn[2985] = 0;
decompressedDataIn[2986] = 0;
decompressedDataIn[2987] = 0;
decompressedDataIn[2988] = 0;
decompressedDataIn[2989] = 0;
decompressedDataIn[2990] = 0;
decompressedDataIn[2991] = 0;
decompressedDataIn[2992] = 0;
decompressedDataIn[2993] = 0;
decompressedDataIn[2994] = 0;
decompressedDataIn[2995] = 0;
decompressedDataIn[2996] = 0;
decompressedDataIn[2997] = 0;
decompressedDataIn[2998] = 0;
decompressedDataIn[2999] = 0;
decompressedDataIn[3000] = 0;
decompressedDataIn[3001] = 0;
decompressedDataIn[3002] = 0;
decompressedDataIn[3003] = 0;
decompressedDataIn[3004] = 0;
decompressedDataIn[3005] = 0;
decompressedDataIn[3006] = 0;
decompressedDataIn[3007] = 0;
decompressedDataIn[3008] = 0;
decompressedDataIn[3009] = 0;
decompressedDataIn[3010] = 0;
decompressedDataIn[3011] = 0;
decompressedDataIn[3012] = 0;
decompressedDataIn[3013] = 0;
decompressedDataIn[3014] = 0;
decompressedDataIn[3015] = 0;
decompressedDataIn[3016] = 0;
decompressedDataIn[3017] = 0;
decompressedDataIn[3018] = 0;
decompressedDataIn[3019] = 0;
decompressedDataIn[3020] = 0;
decompressedDataIn[3021] = 0;
decompressedDataIn[3022] = 0;
decompressedDataIn[3023] = 0;
decompressedDataIn[3024] = 0;
decompressedDataIn[3025] = 0;
decompressedDataIn[3026] = 0;
decompressedDataIn[3027] = 0;
decompressedDataIn[3028] = 0;
decompressedDataIn[3029] = 0;
decompressedDataIn[3030] = 0;
decompressedDataIn[3031] = 0;
decompressedDataIn[3032] = 0;
decompressedDataIn[3033] = 0;
decompressedDataIn[3034] = 0;
decompressedDataIn[3035] = 0;
decompressedDataIn[3036] = 0;
decompressedDataIn[3037] = 0;
decompressedDataIn[3038] = 0;
decompressedDataIn[3039] = 0;
decompressedDataIn[3040] = 0;
decompressedDataIn[3041] = 0;
decompressedDataIn[3042] = 0;
decompressedDataIn[3043] = 0;
decompressedDataIn[3044] = 0;
decompressedDataIn[3045] = 0;
decompressedDataIn[3046] = 0;
decompressedDataIn[3047] = 0;
decompressedDataIn[3048] = 0;
decompressedDataIn[3049] = 0;
decompressedDataIn[3050] = 0;
decompressedDataIn[3051] = 0;
decompressedDataIn[3052] = 0;
decompressedDataIn[3053] = 0;
decompressedDataIn[3054] = 0;
decompressedDataIn[3055] = 0;
decompressedDataIn[3056] = 0;
decompressedDataIn[3057] = 0;
decompressedDataIn[3058] = 0;
decompressedDataIn[3059] = 0;
decompressedDataIn[3060] = 0;
decompressedDataIn[3061] = 0;
decompressedDataIn[3062] = 0;
decompressedDataIn[3063] = 0;
decompressedDataIn[3064] = 0;
decompressedDataIn[3065] = 0;
decompressedDataIn[3066] = 0;
decompressedDataIn[3067] = 0;
decompressedDataIn[3068] = 0;
decompressedDataIn[3069] = 0;
decompressedDataIn[3070] = 0;
decompressedDataIn[3071] = 0;
decompressedDataIn[3072] = 0;
decompressedDataIn[3073] = 0;
decompressedDataIn[3074] = 0;
decompressedDataIn[3075] = 0;
decompressedDataIn[3076] = 0;
decompressedDataIn[3077] = 0;
decompressedDataIn[3078] = 0;
decompressedDataIn[3079] = 0;
decompressedDataIn[3080] = 0;
decompressedDataIn[3081] = 0;
decompressedDataIn[3082] = 0;
decompressedDataIn[3083] = 0;
decompressedDataIn[3084] = 0;
decompressedDataIn[3085] = 0;
decompressedDataIn[3086] = 0;
decompressedDataIn[3087] = 0;
decompressedDataIn[3088] = 0;
decompressedDataIn[3089] = 0;
decompressedDataIn[3090] = 0;
decompressedDataIn[3091] = 0;
decompressedDataIn[3092] = 0;
decompressedDataIn[3093] = 0;
decompressedDataIn[3094] = 0;
decompressedDataIn[3095] = 0;
decompressedDataIn[3096] = 0;
decompressedDataIn[3097] = 0;
decompressedDataIn[3098] = 0;
decompressedDataIn[3099] = 0;
decompressedDataIn[3100] = 0;
decompressedDataIn[3101] = 0;
decompressedDataIn[3102] = 0;
decompressedDataIn[3103] = 0;
decompressedDataIn[3104] = 0;
decompressedDataIn[3105] = 0;
decompressedDataIn[3106] = 0;
decompressedDataIn[3107] = 0;
decompressedDataIn[3108] = 0;
decompressedDataIn[3109] = 0;
decompressedDataIn[3110] = 0;
decompressedDataIn[3111] = 0;
decompressedDataIn[3112] = 0;
decompressedDataIn[3113] = 0;
decompressedDataIn[3114] = 0;
decompressedDataIn[3115] = 0;
decompressedDataIn[3116] = 0;
decompressedDataIn[3117] = 0;
decompressedDataIn[3118] = 0;
decompressedDataIn[3119] = 0;
decompressedDataIn[3120] = 0;
decompressedDataIn[3121] = 0;
decompressedDataIn[3122] = 0;
decompressedDataIn[3123] = 0;
decompressedDataIn[3124] = 0;
decompressedDataIn[3125] = 0;
decompressedDataIn[3126] = 0;
decompressedDataIn[3127] = 0;
decompressedDataIn[3128] = 0;
decompressedDataIn[3129] = 0;
decompressedDataIn[3130] = 0;
decompressedDataIn[3131] = 0;
decompressedDataIn[3132] = 0;
decompressedDataIn[3133] = 0;
decompressedDataIn[3134] = 0;
decompressedDataIn[3135] = 0;
decompressedDataIn[3136] = 0;
decompressedDataIn[3137] = 0;
decompressedDataIn[3138] = 0;
decompressedDataIn[3139] = 0;
decompressedDataIn[3140] = 0;
decompressedDataIn[3141] = 0;
decompressedDataIn[3142] = 0;
decompressedDataIn[3143] = 0;
decompressedDataIn[3144] = 0;
decompressedDataIn[3145] = 0;
decompressedDataIn[3146] = 0;
decompressedDataIn[3147] = 0;
decompressedDataIn[3148] = 0;
decompressedDataIn[3149] = 0;
decompressedDataIn[3150] = 0;
decompressedDataIn[3151] = 0;
decompressedDataIn[3152] = 0;
decompressedDataIn[3153] = 0;
decompressedDataIn[3154] = 0;
decompressedDataIn[3155] = 0;
decompressedDataIn[3156] = 0;
decompressedDataIn[3157] = 0;
decompressedDataIn[3158] = 0;
decompressedDataIn[3159] = 0;
decompressedDataIn[3160] = 0;
decompressedDataIn[3161] = 0;
decompressedDataIn[3162] = 0;
decompressedDataIn[3163] = 0;
decompressedDataIn[3164] = 0;
decompressedDataIn[3165] = 0;
decompressedDataIn[3166] = 0;
decompressedDataIn[3167] = 0;
decompressedDataIn[3168] = 0;
decompressedDataIn[3169] = 0;
decompressedDataIn[3170] = 0;
decompressedDataIn[3171] = 0;
decompressedDataIn[3172] = 0;
decompressedDataIn[3173] = 0;
decompressedDataIn[3174] = 0;
decompressedDataIn[3175] = 0;
decompressedDataIn[3176] = 0;
decompressedDataIn[3177] = 0;
decompressedDataIn[3178] = 0;
decompressedDataIn[3179] = 0;
decompressedDataIn[3180] = 0;
decompressedDataIn[3181] = 0;
decompressedDataIn[3182] = 0;
decompressedDataIn[3183] = 0;
decompressedDataIn[3184] = 0;
decompressedDataIn[3185] = 0;
decompressedDataIn[3186] = 0;
decompressedDataIn[3187] = 0;
decompressedDataIn[3188] = 0;
decompressedDataIn[3189] = 0;
decompressedDataIn[3190] = 0;
decompressedDataIn[3191] = 0;
decompressedDataIn[3192] = 0;
decompressedDataIn[3193] = 0;
decompressedDataIn[3194] = 0;
decompressedDataIn[3195] = 0;
decompressedDataIn[3196] = 0;
decompressedDataIn[3197] = 0;
decompressedDataIn[3198] = 0;
decompressedDataIn[3199] = 0;
decompressedDataIn[3200] = 0;
decompressedDataIn[3201] = 0;
decompressedDataIn[3202] = 0;
decompressedDataIn[3203] = 0;
decompressedDataIn[3204] = 0;
decompressedDataIn[3205] = 0;
decompressedDataIn[3206] = 0;
decompressedDataIn[3207] = 0;
decompressedDataIn[3208] = 0;
decompressedDataIn[3209] = 0;
decompressedDataIn[3210] = 0;
decompressedDataIn[3211] = 0;
decompressedDataIn[3212] = 0;
decompressedDataIn[3213] = 0;
decompressedDataIn[3214] = 0;
decompressedDataIn[3215] = 0;
decompressedDataIn[3216] = 0;
decompressedDataIn[3217] = 0;
decompressedDataIn[3218] = 0;
decompressedDataIn[3219] = 0;
decompressedDataIn[3220] = 0;
decompressedDataIn[3221] = 0;
decompressedDataIn[3222] = 0;
decompressedDataIn[3223] = 0;
decompressedDataIn[3224] = 0;
decompressedDataIn[3225] = 0;
decompressedDataIn[3226] = 0;
decompressedDataIn[3227] = 0;
decompressedDataIn[3228] = 0;
decompressedDataIn[3229] = 0;
decompressedDataIn[3230] = 0;
decompressedDataIn[3231] = 0;
decompressedDataIn[3232] = 0;
decompressedDataIn[3233] = 0;
decompressedDataIn[3234] = 0;
decompressedDataIn[3235] = 0;
decompressedDataIn[3236] = 0;
decompressedDataIn[3237] = 0;
decompressedDataIn[3238] = 0;
decompressedDataIn[3239] = 0;
decompressedDataIn[3240] = 0;
decompressedDataIn[3241] = 0;
decompressedDataIn[3242] = 0;
decompressedDataIn[3243] = 0;
decompressedDataIn[3244] = 0;
decompressedDataIn[3245] = 0;
decompressedDataIn[3246] = 0;
decompressedDataIn[3247] = 0;
decompressedDataIn[3248] = 0;
decompressedDataIn[3249] = 0;
decompressedDataIn[3250] = 0;
decompressedDataIn[3251] = 0;
decompressedDataIn[3252] = 0;
decompressedDataIn[3253] = 0;
decompressedDataIn[3254] = 0;
decompressedDataIn[3255] = 0;
decompressedDataIn[3256] = 0;
decompressedDataIn[3257] = 0;
decompressedDataIn[3258] = 0;
decompressedDataIn[3259] = 0;
decompressedDataIn[3260] = 0;
decompressedDataIn[3261] = 0;
decompressedDataIn[3262] = 0;
decompressedDataIn[3263] = 0;
decompressedDataIn[3264] = 0;
decompressedDataIn[3265] = 0;
decompressedDataIn[3266] = 0;
decompressedDataIn[3267] = 0;
decompressedDataIn[3268] = 0;
decompressedDataIn[3269] = 0;
decompressedDataIn[3270] = 0;
decompressedDataIn[3271] = 0;
decompressedDataIn[3272] = 0;
decompressedDataIn[3273] = 0;
decompressedDataIn[3274] = 0;
decompressedDataIn[3275] = 0;
decompressedDataIn[3276] = 0;
decompressedDataIn[3277] = 0;
decompressedDataIn[3278] = 0;
decompressedDataIn[3279] = 0;
decompressedDataIn[3280] = 0;
decompressedDataIn[3281] = 0;
decompressedDataIn[3282] = 0;
decompressedDataIn[3283] = 0;
decompressedDataIn[3284] = 0;
decompressedDataIn[3285] = 0;
decompressedDataIn[3286] = 0;
decompressedDataIn[3287] = 0;
decompressedDataIn[3288] = 0;
decompressedDataIn[3289] = 0;
decompressedDataIn[3290] = 0;
decompressedDataIn[3291] = 0;
decompressedDataIn[3292] = 0;
decompressedDataIn[3293] = 0;
decompressedDataIn[3294] = 0;
decompressedDataIn[3295] = 0;
decompressedDataIn[3296] = 0;
decompressedDataIn[3297] = 0;
decompressedDataIn[3298] = 0;
decompressedDataIn[3299] = 0;
decompressedDataIn[3300] = 0;
decompressedDataIn[3301] = 0;
decompressedDataIn[3302] = 0;
decompressedDataIn[3303] = 0;
decompressedDataIn[3304] = 0;
decompressedDataIn[3305] = 0;
decompressedDataIn[3306] = 0;
decompressedDataIn[3307] = 0;
decompressedDataIn[3308] = 0;
decompressedDataIn[3309] = 0;
decompressedDataIn[3310] = 0;
decompressedDataIn[3311] = 0;
decompressedDataIn[3312] = 0;
decompressedDataIn[3313] = 0;
decompressedDataIn[3314] = 0;
decompressedDataIn[3315] = 0;
decompressedDataIn[3316] = 0;
decompressedDataIn[3317] = 0;
decompressedDataIn[3318] = 0;
decompressedDataIn[3319] = 0;
decompressedDataIn[3320] = 0;
decompressedDataIn[3321] = 0;
decompressedDataIn[3322] = 0;
decompressedDataIn[3323] = 0;
decompressedDataIn[3324] = 0;
decompressedDataIn[3325] = 0;
decompressedDataIn[3326] = 0;
decompressedDataIn[3327] = 0;
decompressedDataIn[3328] = 0;
decompressedDataIn[3329] = 0;
decompressedDataIn[3330] = 0;
decompressedDataIn[3331] = 0;
decompressedDataIn[3332] = 0;
decompressedDataIn[3333] = 0;
decompressedDataIn[3334] = 0;
decompressedDataIn[3335] = 0;
decompressedDataIn[3336] = 5;
decompressedDataIn[3337] = 0;
decompressedDataIn[3338] = 0;
decompressedDataIn[3339] = 0;
decompressedDataIn[3340] = 128;
decompressedDataIn[3341] = 0;
decompressedDataIn[3342] = 0;
decompressedDataIn[3343] = 0;
decompressedDataIn[3344] = 73;
decompressedDataIn[3345] = 71;
decompressedDataIn[3346] = 73;
decompressedDataIn[3347] = 83;
decompressedDataIn[3348] = 67;
decompressedDataIn[3349] = 79;
decompressedDataIn[3350] = 82;
decompressedDataIn[3351] = 69;
decompressedDataIn[3352] = 0;
decompressedDataIn[3353] = 0;
decompressedDataIn[3354] = 0;
decompressedDataIn[3355] = 0;
decompressedDataIn[3356] = 19;
decompressedDataIn[3357] = 0;
decompressedDataIn[3358] = 0;
decompressedDataIn[3359] = 0;
decompressedDataIn[3360] = 0;
decompressedDataIn[3361] = 0;
decompressedDataIn[3362] = 0;
decompressedDataIn[3363] = 0;
decompressedDataIn[3364] = 128;
decompressedDataIn[3365] = 0;
decompressedDataIn[3366] = 0;
decompressedDataIn[3367] = 0;
decompressedDataIn[3368] = 0;
decompressedDataIn[3369] = 0;
decompressedDataIn[3370] = 0;
decompressedDataIn[3371] = 0;
decompressedDataIn[3372] = 0;
decompressedDataIn[3373] = 0;
decompressedDataIn[3374] = 0;
decompressedDataIn[3375] = 0;
decompressedDataIn[3376] = 0;
decompressedDataIn[3377] = 0;
decompressedDataIn[3378] = 0;
decompressedDataIn[3379] = 0;
decompressedDataIn[3380] = 0;
decompressedDataIn[3381] = 0;
decompressedDataIn[3382] = 0;
decompressedDataIn[3383] = 0;
decompressedDataIn[3384] = 0;
decompressedDataIn[3385] = 0;
decompressedDataIn[3386] = 0;
decompressedDataIn[3387] = 0;
decompressedDataIn[3388] = 0;
decompressedDataIn[3389] = 0;
decompressedDataIn[3390] = 0;
decompressedDataIn[3391] = 0;
decompressedDataIn[3392] = 0;
decompressedDataIn[3393] = 0;
decompressedDataIn[3394] = 0;
decompressedDataIn[3395] = 0;
decompressedDataIn[3396] = 0;
decompressedDataIn[3397] = 0;
decompressedDataIn[3398] = 0;
decompressedDataIn[3399] = 0;
decompressedDataIn[3400] = 0;
decompressedDataIn[3401] = 0;
decompressedDataIn[3402] = 0;
decompressedDataIn[3403] = 0;
decompressedDataIn[3404] = 0;
decompressedDataIn[3405] = 0;
decompressedDataIn[3406] = 0;
decompressedDataIn[3407] = 0;
decompressedDataIn[3408] = 0;
decompressedDataIn[3409] = 0;
decompressedDataIn[3410] = 0;
decompressedDataIn[3411] = 0;
decompressedDataIn[3412] = 0;
decompressedDataIn[3413] = 0;
decompressedDataIn[3414] = 0;
decompressedDataIn[3415] = 0;
decompressedDataIn[3416] = 0;
decompressedDataIn[3417] = 0;
decompressedDataIn[3418] = 0;
decompressedDataIn[3419] = 0;
decompressedDataIn[3420] = 0;
decompressedDataIn[3421] = 0;
decompressedDataIn[3422] = 0;
decompressedDataIn[3423] = 0;
decompressedDataIn[3424] = 0;
decompressedDataIn[3425] = 0;
decompressedDataIn[3426] = 0;
decompressedDataIn[3427] = 0;
decompressedDataIn[3428] = 0;
decompressedDataIn[3429] = 0;
decompressedDataIn[3430] = 0;
decompressedDataIn[3431] = 0;
decompressedDataIn[3432] = 0;
decompressedDataIn[3433] = 0;
decompressedDataIn[3434] = 0;
decompressedDataIn[3435] = 0;
decompressedDataIn[3436] = 0;
decompressedDataIn[3437] = 0;
decompressedDataIn[3438] = 0;
decompressedDataIn[3439] = 0;
decompressedDataIn[3440] = 0;
decompressedDataIn[3441] = 0;
decompressedDataIn[3442] = 0;
decompressedDataIn[3443] = 0;
decompressedDataIn[3444] = 0;
decompressedDataIn[3445] = 0;
decompressedDataIn[3446] = 0;
decompressedDataIn[3447] = 0;
decompressedDataIn[3448] = 0;
decompressedDataIn[3449] = 0;
decompressedDataIn[3450] = 0;
decompressedDataIn[3451] = 0;
decompressedDataIn[3452] = 0;
decompressedDataIn[3453] = 0;
decompressedDataIn[3454] = 0;
decompressedDataIn[3455] = 0;
decompressedDataIn[3456] = 0;
decompressedDataIn[3457] = 0;
decompressedDataIn[3458] = 0;
decompressedDataIn[3459] = 0;
decompressedDataIn[3460] = 0;
decompressedDataIn[3461] = 0;
decompressedDataIn[3462] = 0;
decompressedDataIn[3463] = 0;
decompressedDataIn[3464] = 0;
decompressedDataIn[3465] = 0;
decompressedDataIn[3466] = 0;
decompressedDataIn[3467] = 0;
decompressedDataIn[3468] = 0;
decompressedDataIn[3469] = 0;
decompressedDataIn[3470] = 0;
decompressedDataIn[3471] = 0;
decompressedDataIn[3472] = 0;
decompressedDataIn[3473] = 0;
decompressedDataIn[3474] = 0;
decompressedDataIn[3475] = 0;
decompressedDataIn[3476] = 0;
decompressedDataIn[3477] = 0;
decompressedDataIn[3478] = 0;
decompressedDataIn[3479] = 0;
decompressedDataIn[3480] = 0;
decompressedDataIn[3481] = 0;
decompressedDataIn[3482] = 0;
decompressedDataIn[3483] = 0;
decompressedDataIn[3484] = 5;
decompressedDataIn[3485] = 0;
decompressedDataIn[3486] = 0;
decompressedDataIn[3487] = 0;
decompressedDataIn[3488] = 64;
decompressedDataIn[3489] = 1;
decompressedDataIn[3490] = 0;
decompressedDataIn[3491] = 0;
decompressedDataIn[3492] = 6;
decompressedDataIn[3493] = 0;
decompressedDataIn[3494] = 0;
decompressedDataIn[3495] = 0;
decompressedDataIn[3496] = 67;
decompressedDataIn[3497] = 79;
decompressedDataIn[3498] = 82;
decompressedDataIn[3499] = 69;
decompressedDataIn[3500] = 0;
decompressedDataIn[3501] = 0;
decompressedDataIn[3502] = 0;
decompressedDataIn[3503] = 0;
decompressedDataIn[3504] = 33;
decompressedDataIn[3505] = 0;
decompressedDataIn[3506] = 0;
decompressedDataIn[3507] = 0;
decompressedDataIn[3508] = 0;
decompressedDataIn[3509] = 0;
decompressedDataIn[3510] = 0;
decompressedDataIn[3511] = 0;
decompressedDataIn[3512] = 0;
decompressedDataIn[3513] = 64;
decompressedDataIn[3514] = 94;
decompressedDataIn[3515] = 67;
decompressedDataIn[3516] = 255;
decompressedDataIn[3517] = 127;
decompressedDataIn[3518] = 0;
decompressedDataIn[3519] = 0;
decompressedDataIn[3520] = 16;
decompressedDataIn[3521] = 0;
decompressedDataIn[3522] = 0;
decompressedDataIn[3523] = 0;
decompressedDataIn[3524] = 0;
decompressedDataIn[3525] = 0;
decompressedDataIn[3526] = 0;
decompressedDataIn[3527] = 0;
decompressedDataIn[3528] = 255;
decompressedDataIn[3529] = 251;
decompressedDataIn[3530] = 235;
decompressedDataIn[3531] = 191;
decompressedDataIn[3532] = 0;
decompressedDataIn[3533] = 0;
decompressedDataIn[3534] = 0;
decompressedDataIn[3535] = 0;
decompressedDataIn[3536] = 6;
decompressedDataIn[3537] = 0;
decompressedDataIn[3538] = 0;
decompressedDataIn[3539] = 0;
decompressedDataIn[3540] = 0;
decompressedDataIn[3541] = 0;
decompressedDataIn[3542] = 0;
decompressedDataIn[3543] = 0;
decompressedDataIn[3544] = 0;
decompressedDataIn[3545] = 16;
decompressedDataIn[3546] = 0;
decompressedDataIn[3547] = 0;
decompressedDataIn[3548] = 0;
decompressedDataIn[3549] = 0;
decompressedDataIn[3550] = 0;
decompressedDataIn[3551] = 0;
decompressedDataIn[3552] = 17;
decompressedDataIn[3553] = 0;
decompressedDataIn[3554] = 0;
decompressedDataIn[3555] = 0;
decompressedDataIn[3556] = 0;
decompressedDataIn[3557] = 0;
decompressedDataIn[3558] = 0;
decompressedDataIn[3559] = 0;
decompressedDataIn[3560] = 100;
decompressedDataIn[3561] = 0;
decompressedDataIn[3562] = 0;
decompressedDataIn[3563] = 0;
decompressedDataIn[3564] = 0;
decompressedDataIn[3565] = 0;
decompressedDataIn[3566] = 0;
decompressedDataIn[3567] = 0;
decompressedDataIn[3568] = 3;
decompressedDataIn[3569] = 0;
decompressedDataIn[3570] = 0;
decompressedDataIn[3571] = 0;
decompressedDataIn[3572] = 0;
decompressedDataIn[3573] = 0;
decompressedDataIn[3574] = 0;
decompressedDataIn[3575] = 0;
decompressedDataIn[3576] = 64;
decompressedDataIn[3577] = 0;
decompressedDataIn[3578] = 171;
decompressedDataIn[3579] = 213;
decompressedDataIn[3580] = 109;
decompressedDataIn[3581] = 85;
decompressedDataIn[3582] = 0;
decompressedDataIn[3583] = 0;
decompressedDataIn[3584] = 4;
decompressedDataIn[3585] = 0;
decompressedDataIn[3586] = 0;
decompressedDataIn[3587] = 0;
decompressedDataIn[3588] = 0;
decompressedDataIn[3589] = 0;
decompressedDataIn[3590] = 0;
decompressedDataIn[3591] = 0;
decompressedDataIn[3592] = 56;
decompressedDataIn[3593] = 0;
decompressedDataIn[3594] = 0;
decompressedDataIn[3595] = 0;
decompressedDataIn[3596] = 0;
decompressedDataIn[3597] = 0;
decompressedDataIn[3598] = 0;
decompressedDataIn[3599] = 0;
decompressedDataIn[3600] = 5;
decompressedDataIn[3601] = 0;
decompressedDataIn[3602] = 0;
decompressedDataIn[3603] = 0;
decompressedDataIn[3604] = 0;
decompressedDataIn[3605] = 0;
decompressedDataIn[3606] = 0;
decompressedDataIn[3607] = 0;
decompressedDataIn[3608] = 9;
decompressedDataIn[3609] = 0;
decompressedDataIn[3610] = 0;
decompressedDataIn[3611] = 0;
decompressedDataIn[3612] = 0;
decompressedDataIn[3613] = 0;
decompressedDataIn[3614] = 0;
decompressedDataIn[3615] = 0;
decompressedDataIn[3616] = 7;
decompressedDataIn[3617] = 0;
decompressedDataIn[3618] = 0;
decompressedDataIn[3619] = 0;
decompressedDataIn[3620] = 0;
decompressedDataIn[3621] = 0;
decompressedDataIn[3622] = 0;
decompressedDataIn[3623] = 0;
decompressedDataIn[3624] = 0;
decompressedDataIn[3625] = 32;
decompressedDataIn[3626] = 146;
decompressedDataIn[3627] = 247;
decompressedDataIn[3628] = 217;
decompressedDataIn[3629] = 127;
decompressedDataIn[3630] = 0;
decompressedDataIn[3631] = 0;
decompressedDataIn[3632] = 8;
decompressedDataIn[3633] = 0;
decompressedDataIn[3634] = 0;
decompressedDataIn[3635] = 0;
decompressedDataIn[3636] = 0;
decompressedDataIn[3637] = 0;
decompressedDataIn[3638] = 0;
decompressedDataIn[3639] = 0;
decompressedDataIn[3640] = 0;
decompressedDataIn[3641] = 0;
decompressedDataIn[3642] = 0;
decompressedDataIn[3643] = 0;
decompressedDataIn[3644] = 0;
decompressedDataIn[3645] = 0;
decompressedDataIn[3646] = 0;
decompressedDataIn[3647] = 0;
decompressedDataIn[3648] = 9;
decompressedDataIn[3649] = 0;
decompressedDataIn[3650] = 0;
decompressedDataIn[3651] = 0;
decompressedDataIn[3652] = 0;
decompressedDataIn[3653] = 0;
decompressedDataIn[3654] = 0;
decompressedDataIn[3655] = 0;
decompressedDataIn[3656] = 176;
decompressedDataIn[3657] = 10;
decompressedDataIn[3658] = 171;
decompressedDataIn[3659] = 213;
decompressedDataIn[3660] = 109;
decompressedDataIn[3661] = 85;
decompressedDataIn[3662] = 0;
decompressedDataIn[3663] = 0;
decompressedDataIn[3664] = 11;
decompressedDataIn[3665] = 0;
decompressedDataIn[3666] = 0;
decompressedDataIn[3667] = 0;
decompressedDataIn[3668] = 0;
decompressedDataIn[3669] = 0;
decompressedDataIn[3670] = 0;
decompressedDataIn[3671] = 0;
decompressedDataIn[3672] = 0;
decompressedDataIn[3673] = 0;
decompressedDataIn[3674] = 0;
decompressedDataIn[3675] = 0;
decompressedDataIn[3676] = 0;
decompressedDataIn[3677] = 0;
decompressedDataIn[3678] = 0;
decompressedDataIn[3679] = 0;
decompressedDataIn[3680] = 12;
decompressedDataIn[3681] = 0;
decompressedDataIn[3682] = 0;
decompressedDataIn[3683] = 0;
decompressedDataIn[3684] = 0;
decompressedDataIn[3685] = 0;
decompressedDataIn[3686] = 0;
decompressedDataIn[3687] = 0;
decompressedDataIn[3688] = 0;
decompressedDataIn[3689] = 0;
decompressedDataIn[3690] = 0;
decompressedDataIn[3691] = 0;
decompressedDataIn[3692] = 0;
decompressedDataIn[3693] = 0;
decompressedDataIn[3694] = 0;
decompressedDataIn[3695] = 0;
decompressedDataIn[3696] = 13;
decompressedDataIn[3697] = 0;
decompressedDataIn[3698] = 0;
decompressedDataIn[3699] = 0;
decompressedDataIn[3700] = 0;
decompressedDataIn[3701] = 0;
decompressedDataIn[3702] = 0;
decompressedDataIn[3703] = 0;
decompressedDataIn[3704] = 0;
decompressedDataIn[3705] = 0;
decompressedDataIn[3706] = 0;
decompressedDataIn[3707] = 0;
decompressedDataIn[3708] = 0;
decompressedDataIn[3709] = 0;
decompressedDataIn[3710] = 0;
decompressedDataIn[3711] = 0;
decompressedDataIn[3712] = 14;
decompressedDataIn[3713] = 0;
decompressedDataIn[3714] = 0;
decompressedDataIn[3715] = 0;
decompressedDataIn[3716] = 0;
decompressedDataIn[3717] = 0;
decompressedDataIn[3718] = 0;
decompressedDataIn[3719] = 0;
decompressedDataIn[3720] = 0;
decompressedDataIn[3721] = 0;
decompressedDataIn[3722] = 0;
decompressedDataIn[3723] = 0;
decompressedDataIn[3724] = 0;
decompressedDataIn[3725] = 0;
decompressedDataIn[3726] = 0;
decompressedDataIn[3727] = 0;
decompressedDataIn[3728] = 23;
decompressedDataIn[3729] = 0;
decompressedDataIn[3730] = 0;
decompressedDataIn[3731] = 0;
decompressedDataIn[3732] = 0;
decompressedDataIn[3733] = 0;
decompressedDataIn[3734] = 0;
decompressedDataIn[3735] = 0;
decompressedDataIn[3736] = 0;
decompressedDataIn[3737] = 0;
decompressedDataIn[3738] = 0;
decompressedDataIn[3739] = 0;
decompressedDataIn[3740] = 0;
decompressedDataIn[3741] = 0;
decompressedDataIn[3742] = 0;
decompressedDataIn[3743] = 0;
decompressedDataIn[3744] = 25;
decompressedDataIn[3745] = 0;
decompressedDataIn[3746] = 0;
decompressedDataIn[3747] = 0;
decompressedDataIn[3748] = 0;
decompressedDataIn[3749] = 0;
decompressedDataIn[3750] = 0;
decompressedDataIn[3751] = 0;
decompressedDataIn[3752] = 249;
decompressedDataIn[3753] = 117;
decompressedDataIn[3754] = 67;
decompressedDataIn[3755] = 67;
decompressedDataIn[3756] = 255;
decompressedDataIn[3757] = 127;
decompressedDataIn[3758] = 0;
decompressedDataIn[3759] = 0;
decompressedDataIn[3760] = 26;
decompressedDataIn[3761] = 0;
decompressedDataIn[3762] = 0;
decompressedDataIn[3763] = 0;
decompressedDataIn[3764] = 0;
decompressedDataIn[3765] = 0;
decompressedDataIn[3766] = 0;
decompressedDataIn[3767] = 0;
decompressedDataIn[3768] = 0;
decompressedDataIn[3769] = 0;
decompressedDataIn[3770] = 0;
decompressedDataIn[3771] = 0;
decompressedDataIn[3772] = 0;
decompressedDataIn[3773] = 0;
decompressedDataIn[3774] = 0;
decompressedDataIn[3775] = 0;
decompressedDataIn[3776] = 31;
decompressedDataIn[3777] = 0;
decompressedDataIn[3778] = 0;
decompressedDataIn[3779] = 0;
decompressedDataIn[3780] = 0;
decompressedDataIn[3781] = 0;
decompressedDataIn[3782] = 0;
decompressedDataIn[3783] = 0;
decompressedDataIn[3784] = 136;
decompressedDataIn[3785] = 143;
decompressedDataIn[3786] = 67;
decompressedDataIn[3787] = 67;
decompressedDataIn[3788] = 255;
decompressedDataIn[3789] = 127;
decompressedDataIn[3790] = 0;
decompressedDataIn[3791] = 0;
decompressedDataIn[3792] = 15;
decompressedDataIn[3793] = 0;
decompressedDataIn[3794] = 0;
decompressedDataIn[3795] = 0;
decompressedDataIn[3796] = 0;
decompressedDataIn[3797] = 0;
decompressedDataIn[3798] = 0;
decompressedDataIn[3799] = 0;
decompressedDataIn[3800] = 9;
decompressedDataIn[3801] = 118;
decompressedDataIn[3802] = 67;
decompressedDataIn[3803] = 67;
decompressedDataIn[3804] = 255;
decompressedDataIn[3805] = 127;
decompressedDataIn[3806] = 0;
decompressedDataIn[3807] = 0;
decompressedDataIn[3808] = 0;
decompressedDataIn[3809] = 0;
decompressedDataIn[3810] = 0;
decompressedDataIn[3811] = 0;
decompressedDataIn[3812] = 0;
decompressedDataIn[3813] = 0;
decompressedDataIn[3814] = 0;
decompressedDataIn[3815] = 0;
decompressedDataIn[3816] = 0;
decompressedDataIn[3817] = 0;
decompressedDataIn[3818] = 0;
decompressedDataIn[3819] = 0;
decompressedDataIn[3820] = 0;
decompressedDataIn[3821] = 0;
decompressedDataIn[3822] = 0;
decompressedDataIn[3823] = 0;
decompressedDataIn[3824] = 5;
decompressedDataIn[3825] = 0;
decompressedDataIn[3826] = 0;
decompressedDataIn[3827] = 0;
decompressedDataIn[3828] = 0;
decompressedDataIn[3829] = 3;
decompressedDataIn[3830] = 0;
decompressedDataIn[3831] = 0;
decompressedDataIn[3832] = 69;
decompressedDataIn[3833] = 76;
decompressedDataIn[3834] = 73;
decompressedDataIn[3835] = 70;
decompressedDataIn[3836] = 67;
decompressedDataIn[3837] = 79;
decompressedDataIn[3838] = 82;
decompressedDataIn[3839] = 69;
decompressedDataIn[3840] = 0;
decompressedDataIn[3841] = 0;
decompressedDataIn[3842] = 0;
decompressedDataIn[3843] = 0;
decompressedDataIn[3844] = 10;
decompressedDataIn[3845] = 0;
decompressedDataIn[3846] = 0;
decompressedDataIn[3847] = 0;
decompressedDataIn[3848] = 0;
decompressedDataIn[3849] = 0;
decompressedDataIn[3850] = 0;
decompressedDataIn[3851] = 0;
decompressedDataIn[3852] = 1;
decompressedDataIn[3853] = 0;
decompressedDataIn[3854] = 0;
decompressedDataIn[3855] = 0;
decompressedDataIn[3856] = 0;
decompressedDataIn[3857] = 0;
decompressedDataIn[3858] = 0;
decompressedDataIn[3859] = 0;
decompressedDataIn[3860] = 0;
decompressedDataIn[3861] = 32;
decompressedDataIn[3862] = 203;
decompressedDataIn[3863] = 213;
decompressedDataIn[3864] = 109;
decompressedDataIn[3865] = 85;
decompressedDataIn[3866] = 0;
decompressedDataIn[3867] = 0;
decompressedDataIn[3868] = 0;
decompressedDataIn[3869] = 48;
decompressedDataIn[3870] = 203;
decompressedDataIn[3871] = 213;
decompressedDataIn[3872] = 109;
decompressedDataIn[3873] = 85;
decompressedDataIn[3874] = 0;
decompressedDataIn[3875] = 0;
decompressedDataIn[3876] = 0;
decompressedDataIn[3877] = 32;
decompressedDataIn[3878] = 0;
decompressedDataIn[3879] = 0;
decompressedDataIn[3880] = 0;
decompressedDataIn[3881] = 0;
decompressedDataIn[3882] = 0;
decompressedDataIn[3883] = 0;
decompressedDataIn[3884] = 0;
decompressedDataIn[3885] = 48;
decompressedDataIn[3886] = 203;
decompressedDataIn[3887] = 213;
decompressedDataIn[3888] = 109;
decompressedDataIn[3889] = 85;
decompressedDataIn[3890] = 0;
decompressedDataIn[3891] = 0;
decompressedDataIn[3892] = 0;
decompressedDataIn[3893] = 64;
decompressedDataIn[3894] = 203;
decompressedDataIn[3895] = 213;
decompressedDataIn[3896] = 109;
decompressedDataIn[3897] = 85;
decompressedDataIn[3898] = 0;
decompressedDataIn[3899] = 0;
decompressedDataIn[3900] = 0;
decompressedDataIn[3901] = 48;
decompressedDataIn[3902] = 0;
decompressedDataIn[3903] = 0;
decompressedDataIn[3904] = 0;
decompressedDataIn[3905] = 0;
decompressedDataIn[3906] = 0;
decompressedDataIn[3907] = 0;
decompressedDataIn[3908] = 0;
decompressedDataIn[3909] = 176;
decompressedDataIn[3910] = 53;
decompressedDataIn[3911] = 247;
decompressedDataIn[3912] = 217;
decompressedDataIn[3913] = 127;
decompressedDataIn[3914] = 0;
decompressedDataIn[3915] = 0;
decompressedDataIn[3916] = 0;
decompressedDataIn[3917] = 240;
decompressedDataIn[3918] = 53;
decompressedDataIn[3919] = 247;
decompressedDataIn[3920] = 217;
decompressedDataIn[3921] = 127;
decompressedDataIn[3922] = 0;
decompressedDataIn[3923] = 0;
decompressedDataIn[3924] = 0;
decompressedDataIn[3925] = 112;
decompressedDataIn[3926] = 30;
decompressedDataIn[3927] = 0;
decompressedDataIn[3928] = 0;
decompressedDataIn[3929] = 0;
decompressedDataIn[3930] = 0;
decompressedDataIn[3931] = 0;
decompressedDataIn[3932] = 0;
decompressedDataIn[3933] = 240;
decompressedDataIn[3934] = 53;
decompressedDataIn[3935] = 247;
decompressedDataIn[3936] = 217;
decompressedDataIn[3937] = 127;
decompressedDataIn[3938] = 0;
decompressedDataIn[3939] = 0;
decompressedDataIn[3940] = 0;
decompressedDataIn[3941] = 16;
decompressedDataIn[3942] = 54;
decompressedDataIn[3943] = 247;
decompressedDataIn[3944] = 217;
decompressedDataIn[3945] = 127;
decompressedDataIn[3946] = 0;
decompressedDataIn[3947] = 0;
decompressedDataIn[3948] = 0;
decompressedDataIn[3949] = 176;
decompressedDataIn[3950] = 30;
decompressedDataIn[3951] = 0;
decompressedDataIn[3952] = 0;
decompressedDataIn[3953] = 0;
decompressedDataIn[3954] = 0;
decompressedDataIn[3955] = 0;
decompressedDataIn[3956] = 0;
decompressedDataIn[3957] = 224;
decompressedDataIn[3958] = 87;
decompressedDataIn[3959] = 247;
decompressedDataIn[3960] = 217;
decompressedDataIn[3961] = 127;
decompressedDataIn[3962] = 0;
decompressedDataIn[3963] = 0;
decompressedDataIn[3964] = 0;
decompressedDataIn[3965] = 240;
decompressedDataIn[3966] = 87;
decompressedDataIn[3967] = 247;
decompressedDataIn[3968] = 217;
decompressedDataIn[3969] = 127;
decompressedDataIn[3970] = 0;
decompressedDataIn[3971] = 0;
decompressedDataIn[3972] = 0;
decompressedDataIn[3973] = 144;
decompressedDataIn[3974] = 1;
decompressedDataIn[3975] = 0;
decompressedDataIn[3976] = 0;
decompressedDataIn[3977] = 0;
decompressedDataIn[3978] = 0;
decompressedDataIn[3979] = 0;
decompressedDataIn[3980] = 0;
decompressedDataIn[3981] = 240;
decompressedDataIn[3982] = 87;
decompressedDataIn[3983] = 247;
decompressedDataIn[3984] = 217;
decompressedDataIn[3985] = 127;
decompressedDataIn[3986] = 0;
decompressedDataIn[3987] = 0;
decompressedDataIn[3988] = 0;
decompressedDataIn[3989] = 0;
decompressedDataIn[3990] = 88;
decompressedDataIn[3991] = 247;
decompressedDataIn[3992] = 217;
decompressedDataIn[3993] = 127;
decompressedDataIn[3994] = 0;
decompressedDataIn[3995] = 0;
decompressedDataIn[3996] = 0;
decompressedDataIn[3997] = 160;
decompressedDataIn[3998] = 1;
decompressedDataIn[3999] = 0;
decompressedDataIn[4000] = 0;
decompressedDataIn[4001] = 0;
decompressedDataIn[4002] = 0;
decompressedDataIn[4003] = 0;
decompressedDataIn[4004] = 0;
decompressedDataIn[4005] = 0;
decompressedDataIn[4006] = 146;
decompressedDataIn[4007] = 247;
decompressedDataIn[4008] = 217;
decompressedDataIn[4009] = 127;
decompressedDataIn[4010] = 0;
decompressedDataIn[4011] = 0;
decompressedDataIn[4012] = 0;
decompressedDataIn[4013] = 16;
decompressedDataIn[4014] = 146;
decompressedDataIn[4015] = 247;
decompressedDataIn[4016] = 217;
decompressedDataIn[4017] = 127;
decompressedDataIn[4018] = 0;
decompressedDataIn[4019] = 0;
decompressedDataIn[4020] = 0;
decompressedDataIn[4021] = 192;
decompressedDataIn[4022] = 25;
decompressedDataIn[4023] = 0;
decompressedDataIn[4024] = 0;
decompressedDataIn[4025] = 0;
decompressedDataIn[4026] = 0;
decompressedDataIn[4027] = 0;
decompressedDataIn[4028] = 0;
decompressedDataIn[4029] = 16;
decompressedDataIn[4030] = 146;
decompressedDataIn[4031] = 247;
decompressedDataIn[4032] = 217;
decompressedDataIn[4033] = 127;
decompressedDataIn[4034] = 0;
decompressedDataIn[4035] = 0;
decompressedDataIn[4036] = 0;
decompressedDataIn[4037] = 32;
decompressedDataIn[4038] = 146;
decompressedDataIn[4039] = 247;
decompressedDataIn[4040] = 217;
decompressedDataIn[4041] = 127;
decompressedDataIn[4042] = 0;
decompressedDataIn[4043] = 0;
decompressedDataIn[4044] = 0;
decompressedDataIn[4045] = 208;
decompressedDataIn[4046] = 25;
decompressedDataIn[4047] = 0;
decompressedDataIn[4048] = 0;
decompressedDataIn[4049] = 0;
decompressedDataIn[4050] = 0;
decompressedDataIn[4051] = 0;
decompressedDataIn[4052] = 0;
decompressedDataIn[4053] = 144;
decompressedDataIn[4054] = 180;
decompressedDataIn[4055] = 247;
decompressedDataIn[4056] = 217;
decompressedDataIn[4057] = 127;
decompressedDataIn[4058] = 0;
decompressedDataIn[4059] = 0;
decompressedDataIn[4060] = 0;
decompressedDataIn[4061] = 160;
decompressedDataIn[4062] = 180;
decompressedDataIn[4063] = 247;
decompressedDataIn[4064] = 217;
decompressedDataIn[4065] = 127;
decompressedDataIn[4066] = 0;
decompressedDataIn[4067] = 0;
decompressedDataIn[4068] = 0;
decompressedDataIn[4069] = 112;
decompressedDataIn[4070] = 2;
decompressedDataIn[4071] = 0;
decompressedDataIn[4072] = 0;
decompressedDataIn[4073] = 0;
decompressedDataIn[4074] = 0;
decompressedDataIn[4075] = 0;
decompressedDataIn[4076] = 0;
decompressedDataIn[4077] = 160;
decompressedDataIn[4078] = 180;
decompressedDataIn[4079] = 247;
decompressedDataIn[4080] = 217;
decompressedDataIn[4081] = 127;
decompressedDataIn[4082] = 0;
decompressedDataIn[4083] = 0;
decompressedDataIn[4084] = 0;
decompressedDataIn[4085] = 176;
decompressedDataIn[4086] = 180;
decompressedDataIn[4087] = 247;
decompressedDataIn[4088] = 217;
decompressedDataIn[4089] = 127;
decompressedDataIn[4090] = 0;
decompressedDataIn[4091] = 0;
decompressedDataIn[4092] = 0;
decompressedDataIn[4093] = 128;
decompressedDataIn[4094] = 2;
decompressedDataIn[4095] = 0;
*/
file = $fopen("testbenchInputFile.txt", "rb");
for(loopCount = 0; loopCount <= desiredLoop; loopCount = loopCount + 1) begin
    r = $fread(decompressedDataIn, file);
end
$fclose(file);
    $display("testinghello");
    #10;
    $display("testinggoodbye");
    clock = 0;
    start = 0;
    #10;
    $display("testing");
    clock = 1;
    #10;
    $display("testing");
    clock = 0;
    start = 1;
    #10;
    $display("testing");
    clock = 1;
    #10;
    $display("testing");
    clock = 0;
    start = 0;
    for(clockCount = 0; clockCount < 100000; clockCount = clockCount + 1)
      begin
    $display("testing%d", clockCount);
        #10;
        clock = 1;
        #10;
        clock = 0;
	if(decompressorFinished && !decompressorFinishedPrevious) begin
		if(inputEqualsOutput) begin
			$display("passed");
		end
		else begin
			$display("failed");
		end
		$finish();
	end
      end
  end

endmodule
