// Wrapper for the toplevel module, which is the combination of the chisel
// implementation for the codeword generator and the compressorOutput

module lzwAndHuffmanWrapper(
         input clock,
         input reset,
         input start,
         input [7:0] dataIn [0:4095],
         output [7:0] dataOut [0:4095],
         output matchBytes [0:4095],
         output [12:0] completeMatch,
         output [12:0] outputBytes,
         output finished,
// These are statistics ports that can easily be disabled and commented out.
	output [10:0] huffmanCharacterDepths [0:16],
	output [3:0] escapeCharacterLength,
	output [5:0] huffmanTreeCharactersUsed,
	output [9:0] dictionaryEntries,
	output [4:0] longestSequenceLength,
	output [12:0] lzUncompressedBytes,
	output [12:0] lzCompressedBytes,
	output [12:0] huffmanCompressedBytes,
       output [13:0] sequenceLengths_0,
       output [13:0] sequenceLengths_1,
       output [13:0] sequenceLengths_2,
       output [13:0] sequenceLengths_3,
       output [13:0] sequenceLengths_4,
       output [13:0] sequenceLengths_5,
       output [13:0] sequenceLengths_6,
       output [13:0] sequenceLengths_7,
       output [13:0] sequenceLengths_8,
       output [13:0] sequenceLengths_9,
       output [13:0] sequenceLengths_10,
       output [13:0] sequenceLengths_11,
       output [13:0] sequenceLengths_12,
       output [13:0] sequenceLengths_13,
       output [13:0] sequenceLengths_14,
       output [13:0] sequenceLengths_15
       );
       wire inValid, inReady, outReady, outValid;

lzwAndHuffman wrapped(
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_0(huffmanCharacterDepths[0]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_1(huffmanCharacterDepths[1]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_2(huffmanCharacterDepths[2]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_3(huffmanCharacterDepths[3]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_4(huffmanCharacterDepths[4]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_5(huffmanCharacterDepths[5]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_6(huffmanCharacterDepths[6]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_7(huffmanCharacterDepths[7]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_8(huffmanCharacterDepths[8]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_9(huffmanCharacterDepths[9]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_10(huffmanCharacterDepths[10]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_11(huffmanCharacterDepths[11]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_12(huffmanCharacterDepths[12]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_13(huffmanCharacterDepths[13]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_14(huffmanCharacterDepths[14]),
.io_compressionStatistics_huffmanStatistics_huffmanCharacterDepths_15(huffmanCharacterDepths[15]),
.io_compressionStatistics_huffmanStatistics_escapeCharacterLength(escapeCharacterLength),
.io_compressionStatistics_huffmanStatistics_huffmanTreeCharactersUsed(huffmanTreeCharactersUsed),
.io_compressionStatistics_lzStatistics_dictionaryEntries(dictionaryEntries),
.io_compressionStatistics_lzStatistics_longestSequenceLength(longestSequenceLength),
.io_compressionStatistics_lzUncompressedBytes(lzUncompressedBytes),
.io_compressionStatistics_lzCompressedBytes(lzCompressedBytes),
.io_compressionStatistics_huffmanCompressedBytes(huffmanCompressedBytes),
.io_compressionStatistics_lzStatistics_sequenceLengths_0(sequenceLengths_0),
.io_compressionStatistics_lzStatistics_sequenceLengths_1(sequenceLengths_1),
.io_compressionStatistics_lzStatistics_sequenceLengths_2(sequenceLengths_2),
.io_compressionStatistics_lzStatistics_sequenceLengths_3(sequenceLengths_3),
.io_compressionStatistics_lzStatistics_sequenceLengths_4(sequenceLengths_4),
.io_compressionStatistics_lzStatistics_sequenceLengths_5(sequenceLengths_5),
.io_compressionStatistics_lzStatistics_sequenceLengths_6(sequenceLengths_6),
.io_compressionStatistics_lzStatistics_sequenceLengths_7(sequenceLengths_7),
.io_compressionStatistics_lzStatistics_sequenceLengths_8(sequenceLengths_8),
.io_compressionStatistics_lzStatistics_sequenceLengths_9(sequenceLengths_9),
.io_compressionStatistics_lzStatistics_sequenceLengths_10(sequenceLengths_10),
.io_compressionStatistics_lzStatistics_sequenceLengths_11(sequenceLengths_11),
.io_compressionStatistics_lzStatistics_sequenceLengths_12(sequenceLengths_12),
.io_compressionStatistics_lzStatistics_sequenceLengths_13(sequenceLengths_13),
.io_compressionStatistics_lzStatistics_sequenceLengths_14(sequenceLengths_14),
.io_compressionStatistics_lzStatistics_sequenceLengths_15(sequenceLengths_15),
.io_start(start),
.clock(clock),
.reset(reset),
.io_parallelIn_0(dataIn[0]),
.io_parallelIn_1(dataIn[1]),
.io_parallelIn_2(dataIn[2]),
.io_parallelIn_3(dataIn[3]),
.io_parallelIn_4(dataIn[4]),
.io_parallelIn_5(dataIn[5]),
.io_parallelIn_6(dataIn[6]),
.io_parallelIn_7(dataIn[7]),
.io_parallelIn_8(dataIn[8]),
.io_parallelIn_9(dataIn[9]),
.io_parallelIn_10(dataIn[10]),
.io_parallelIn_11(dataIn[11]),
.io_parallelIn_12(dataIn[12]),
.io_parallelIn_13(dataIn[13]),
.io_parallelIn_14(dataIn[14]),
.io_parallelIn_15(dataIn[15]),
.io_parallelIn_16(dataIn[16]),
.io_parallelIn_17(dataIn[17]),
.io_parallelIn_18(dataIn[18]),
.io_parallelIn_19(dataIn[19]),
.io_parallelIn_20(dataIn[20]),
.io_parallelIn_21(dataIn[21]),
.io_parallelIn_22(dataIn[22]),
.io_parallelIn_23(dataIn[23]),
.io_parallelIn_24(dataIn[24]),
.io_parallelIn_25(dataIn[25]),
.io_parallelIn_26(dataIn[26]),
.io_parallelIn_27(dataIn[27]),
.io_parallelIn_28(dataIn[28]),
.io_parallelIn_29(dataIn[29]),
.io_parallelIn_30(dataIn[30]),
.io_parallelIn_31(dataIn[31]),
.io_parallelIn_32(dataIn[32]),
.io_parallelIn_33(dataIn[33]),
.io_parallelIn_34(dataIn[34]),
.io_parallelIn_35(dataIn[35]),
.io_parallelIn_36(dataIn[36]),
.io_parallelIn_37(dataIn[37]),
.io_parallelIn_38(dataIn[38]),
.io_parallelIn_39(dataIn[39]),
.io_parallelIn_40(dataIn[40]),
.io_parallelIn_41(dataIn[41]),
.io_parallelIn_42(dataIn[42]),
.io_parallelIn_43(dataIn[43]),
.io_parallelIn_44(dataIn[44]),
.io_parallelIn_45(dataIn[45]),
.io_parallelIn_46(dataIn[46]),
.io_parallelIn_47(dataIn[47]),
.io_parallelIn_48(dataIn[48]),
.io_parallelIn_49(dataIn[49]),
.io_parallelIn_50(dataIn[50]),
.io_parallelIn_51(dataIn[51]),
.io_parallelIn_52(dataIn[52]),
.io_parallelIn_53(dataIn[53]),
.io_parallelIn_54(dataIn[54]),
.io_parallelIn_55(dataIn[55]),
.io_parallelIn_56(dataIn[56]),
.io_parallelIn_57(dataIn[57]),
.io_parallelIn_58(dataIn[58]),
.io_parallelIn_59(dataIn[59]),
.io_parallelIn_60(dataIn[60]),
.io_parallelIn_61(dataIn[61]),
.io_parallelIn_62(dataIn[62]),
.io_parallelIn_63(dataIn[63]),
.io_parallelIn_64(dataIn[64]),
.io_parallelIn_65(dataIn[65]),
.io_parallelIn_66(dataIn[66]),
.io_parallelIn_67(dataIn[67]),
.io_parallelIn_68(dataIn[68]),
.io_parallelIn_69(dataIn[69]),
.io_parallelIn_70(dataIn[70]),
.io_parallelIn_71(dataIn[71]),
.io_parallelIn_72(dataIn[72]),
.io_parallelIn_73(dataIn[73]),
.io_parallelIn_74(dataIn[74]),
.io_parallelIn_75(dataIn[75]),
.io_parallelIn_76(dataIn[76]),
.io_parallelIn_77(dataIn[77]),
.io_parallelIn_78(dataIn[78]),
.io_parallelIn_79(dataIn[79]),
.io_parallelIn_80(dataIn[80]),
.io_parallelIn_81(dataIn[81]),
.io_parallelIn_82(dataIn[82]),
.io_parallelIn_83(dataIn[83]),
.io_parallelIn_84(dataIn[84]),
.io_parallelIn_85(dataIn[85]),
.io_parallelIn_86(dataIn[86]),
.io_parallelIn_87(dataIn[87]),
.io_parallelIn_88(dataIn[88]),
.io_parallelIn_89(dataIn[89]),
.io_parallelIn_90(dataIn[90]),
.io_parallelIn_91(dataIn[91]),
.io_parallelIn_92(dataIn[92]),
.io_parallelIn_93(dataIn[93]),
.io_parallelIn_94(dataIn[94]),
.io_parallelIn_95(dataIn[95]),
.io_parallelIn_96(dataIn[96]),
.io_parallelIn_97(dataIn[97]),
.io_parallelIn_98(dataIn[98]),
.io_parallelIn_99(dataIn[99]),
.io_parallelIn_100(dataIn[100]),
.io_parallelIn_101(dataIn[101]),
.io_parallelIn_102(dataIn[102]),
.io_parallelIn_103(dataIn[103]),
.io_parallelIn_104(dataIn[104]),
.io_parallelIn_105(dataIn[105]),
.io_parallelIn_106(dataIn[106]),
.io_parallelIn_107(dataIn[107]),
.io_parallelIn_108(dataIn[108]),
.io_parallelIn_109(dataIn[109]),
.io_parallelIn_110(dataIn[110]),
.io_parallelIn_111(dataIn[111]),
.io_parallelIn_112(dataIn[112]),
.io_parallelIn_113(dataIn[113]),
.io_parallelIn_114(dataIn[114]),
.io_parallelIn_115(dataIn[115]),
.io_parallelIn_116(dataIn[116]),
.io_parallelIn_117(dataIn[117]),
.io_parallelIn_118(dataIn[118]),
.io_parallelIn_119(dataIn[119]),
.io_parallelIn_120(dataIn[120]),
.io_parallelIn_121(dataIn[121]),
.io_parallelIn_122(dataIn[122]),
.io_parallelIn_123(dataIn[123]),
.io_parallelIn_124(dataIn[124]),
.io_parallelIn_125(dataIn[125]),
.io_parallelIn_126(dataIn[126]),
.io_parallelIn_127(dataIn[127]),
.io_parallelIn_128(dataIn[128]),
.io_parallelIn_129(dataIn[129]),
.io_parallelIn_130(dataIn[130]),
.io_parallelIn_131(dataIn[131]),
.io_parallelIn_132(dataIn[132]),
.io_parallelIn_133(dataIn[133]),
.io_parallelIn_134(dataIn[134]),
.io_parallelIn_135(dataIn[135]),
.io_parallelIn_136(dataIn[136]),
.io_parallelIn_137(dataIn[137]),
.io_parallelIn_138(dataIn[138]),
.io_parallelIn_139(dataIn[139]),
.io_parallelIn_140(dataIn[140]),
.io_parallelIn_141(dataIn[141]),
.io_parallelIn_142(dataIn[142]),
.io_parallelIn_143(dataIn[143]),
.io_parallelIn_144(dataIn[144]),
.io_parallelIn_145(dataIn[145]),
.io_parallelIn_146(dataIn[146]),
.io_parallelIn_147(dataIn[147]),
.io_parallelIn_148(dataIn[148]),
.io_parallelIn_149(dataIn[149]),
.io_parallelIn_150(dataIn[150]),
.io_parallelIn_151(dataIn[151]),
.io_parallelIn_152(dataIn[152]),
.io_parallelIn_153(dataIn[153]),
.io_parallelIn_154(dataIn[154]),
.io_parallelIn_155(dataIn[155]),
.io_parallelIn_156(dataIn[156]),
.io_parallelIn_157(dataIn[157]),
.io_parallelIn_158(dataIn[158]),
.io_parallelIn_159(dataIn[159]),
.io_parallelIn_160(dataIn[160]),
.io_parallelIn_161(dataIn[161]),
.io_parallelIn_162(dataIn[162]),
.io_parallelIn_163(dataIn[163]),
.io_parallelIn_164(dataIn[164]),
.io_parallelIn_165(dataIn[165]),
.io_parallelIn_166(dataIn[166]),
.io_parallelIn_167(dataIn[167]),
.io_parallelIn_168(dataIn[168]),
.io_parallelIn_169(dataIn[169]),
.io_parallelIn_170(dataIn[170]),
.io_parallelIn_171(dataIn[171]),
.io_parallelIn_172(dataIn[172]),
.io_parallelIn_173(dataIn[173]),
.io_parallelIn_174(dataIn[174]),
.io_parallelIn_175(dataIn[175]),
.io_parallelIn_176(dataIn[176]),
.io_parallelIn_177(dataIn[177]),
.io_parallelIn_178(dataIn[178]),
.io_parallelIn_179(dataIn[179]),
.io_parallelIn_180(dataIn[180]),
.io_parallelIn_181(dataIn[181]),
.io_parallelIn_182(dataIn[182]),
.io_parallelIn_183(dataIn[183]),
.io_parallelIn_184(dataIn[184]),
.io_parallelIn_185(dataIn[185]),
.io_parallelIn_186(dataIn[186]),
.io_parallelIn_187(dataIn[187]),
.io_parallelIn_188(dataIn[188]),
.io_parallelIn_189(dataIn[189]),
.io_parallelIn_190(dataIn[190]),
.io_parallelIn_191(dataIn[191]),
.io_parallelIn_192(dataIn[192]),
.io_parallelIn_193(dataIn[193]),
.io_parallelIn_194(dataIn[194]),
.io_parallelIn_195(dataIn[195]),
.io_parallelIn_196(dataIn[196]),
.io_parallelIn_197(dataIn[197]),
.io_parallelIn_198(dataIn[198]),
.io_parallelIn_199(dataIn[199]),
.io_parallelIn_200(dataIn[200]),
.io_parallelIn_201(dataIn[201]),
.io_parallelIn_202(dataIn[202]),
.io_parallelIn_203(dataIn[203]),
.io_parallelIn_204(dataIn[204]),
.io_parallelIn_205(dataIn[205]),
.io_parallelIn_206(dataIn[206]),
.io_parallelIn_207(dataIn[207]),
.io_parallelIn_208(dataIn[208]),
.io_parallelIn_209(dataIn[209]),
.io_parallelIn_210(dataIn[210]),
.io_parallelIn_211(dataIn[211]),
.io_parallelIn_212(dataIn[212]),
.io_parallelIn_213(dataIn[213]),
.io_parallelIn_214(dataIn[214]),
.io_parallelIn_215(dataIn[215]),
.io_parallelIn_216(dataIn[216]),
.io_parallelIn_217(dataIn[217]),
.io_parallelIn_218(dataIn[218]),
.io_parallelIn_219(dataIn[219]),
.io_parallelIn_220(dataIn[220]),
.io_parallelIn_221(dataIn[221]),
.io_parallelIn_222(dataIn[222]),
.io_parallelIn_223(dataIn[223]),
.io_parallelIn_224(dataIn[224]),
.io_parallelIn_225(dataIn[225]),
.io_parallelIn_226(dataIn[226]),
.io_parallelIn_227(dataIn[227]),
.io_parallelIn_228(dataIn[228]),
.io_parallelIn_229(dataIn[229]),
.io_parallelIn_230(dataIn[230]),
.io_parallelIn_231(dataIn[231]),
.io_parallelIn_232(dataIn[232]),
.io_parallelIn_233(dataIn[233]),
.io_parallelIn_234(dataIn[234]),
.io_parallelIn_235(dataIn[235]),
.io_parallelIn_236(dataIn[236]),
.io_parallelIn_237(dataIn[237]),
.io_parallelIn_238(dataIn[238]),
.io_parallelIn_239(dataIn[239]),
.io_parallelIn_240(dataIn[240]),
.io_parallelIn_241(dataIn[241]),
.io_parallelIn_242(dataIn[242]),
.io_parallelIn_243(dataIn[243]),
.io_parallelIn_244(dataIn[244]),
.io_parallelIn_245(dataIn[245]),
.io_parallelIn_246(dataIn[246]),
.io_parallelIn_247(dataIn[247]),
.io_parallelIn_248(dataIn[248]),
.io_parallelIn_249(dataIn[249]),
.io_parallelIn_250(dataIn[250]),
.io_parallelIn_251(dataIn[251]),
.io_parallelIn_252(dataIn[252]),
.io_parallelIn_253(dataIn[253]),
.io_parallelIn_254(dataIn[254]),
.io_parallelIn_255(dataIn[255]),
.io_parallelIn_256(dataIn[256]),
.io_parallelIn_257(dataIn[257]),
.io_parallelIn_258(dataIn[258]),
.io_parallelIn_259(dataIn[259]),
.io_parallelIn_260(dataIn[260]),
.io_parallelIn_261(dataIn[261]),
.io_parallelIn_262(dataIn[262]),
.io_parallelIn_263(dataIn[263]),
.io_parallelIn_264(dataIn[264]),
.io_parallelIn_265(dataIn[265]),
.io_parallelIn_266(dataIn[266]),
.io_parallelIn_267(dataIn[267]),
.io_parallelIn_268(dataIn[268]),
.io_parallelIn_269(dataIn[269]),
.io_parallelIn_270(dataIn[270]),
.io_parallelIn_271(dataIn[271]),
.io_parallelIn_272(dataIn[272]),
.io_parallelIn_273(dataIn[273]),
.io_parallelIn_274(dataIn[274]),
.io_parallelIn_275(dataIn[275]),
.io_parallelIn_276(dataIn[276]),
.io_parallelIn_277(dataIn[277]),
.io_parallelIn_278(dataIn[278]),
.io_parallelIn_279(dataIn[279]),
.io_parallelIn_280(dataIn[280]),
.io_parallelIn_281(dataIn[281]),
.io_parallelIn_282(dataIn[282]),
.io_parallelIn_283(dataIn[283]),
.io_parallelIn_284(dataIn[284]),
.io_parallelIn_285(dataIn[285]),
.io_parallelIn_286(dataIn[286]),
.io_parallelIn_287(dataIn[287]),
.io_parallelIn_288(dataIn[288]),
.io_parallelIn_289(dataIn[289]),
.io_parallelIn_290(dataIn[290]),
.io_parallelIn_291(dataIn[291]),
.io_parallelIn_292(dataIn[292]),
.io_parallelIn_293(dataIn[293]),
.io_parallelIn_294(dataIn[294]),
.io_parallelIn_295(dataIn[295]),
.io_parallelIn_296(dataIn[296]),
.io_parallelIn_297(dataIn[297]),
.io_parallelIn_298(dataIn[298]),
.io_parallelIn_299(dataIn[299]),
.io_parallelIn_300(dataIn[300]),
.io_parallelIn_301(dataIn[301]),
.io_parallelIn_302(dataIn[302]),
.io_parallelIn_303(dataIn[303]),
.io_parallelIn_304(dataIn[304]),
.io_parallelIn_305(dataIn[305]),
.io_parallelIn_306(dataIn[306]),
.io_parallelIn_307(dataIn[307]),
.io_parallelIn_308(dataIn[308]),
.io_parallelIn_309(dataIn[309]),
.io_parallelIn_310(dataIn[310]),
.io_parallelIn_311(dataIn[311]),
.io_parallelIn_312(dataIn[312]),
.io_parallelIn_313(dataIn[313]),
.io_parallelIn_314(dataIn[314]),
.io_parallelIn_315(dataIn[315]),
.io_parallelIn_316(dataIn[316]),
.io_parallelIn_317(dataIn[317]),
.io_parallelIn_318(dataIn[318]),
.io_parallelIn_319(dataIn[319]),
.io_parallelIn_320(dataIn[320]),
.io_parallelIn_321(dataIn[321]),
.io_parallelIn_322(dataIn[322]),
.io_parallelIn_323(dataIn[323]),
.io_parallelIn_324(dataIn[324]),
.io_parallelIn_325(dataIn[325]),
.io_parallelIn_326(dataIn[326]),
.io_parallelIn_327(dataIn[327]),
.io_parallelIn_328(dataIn[328]),
.io_parallelIn_329(dataIn[329]),
.io_parallelIn_330(dataIn[330]),
.io_parallelIn_331(dataIn[331]),
.io_parallelIn_332(dataIn[332]),
.io_parallelIn_333(dataIn[333]),
.io_parallelIn_334(dataIn[334]),
.io_parallelIn_335(dataIn[335]),
.io_parallelIn_336(dataIn[336]),
.io_parallelIn_337(dataIn[337]),
.io_parallelIn_338(dataIn[338]),
.io_parallelIn_339(dataIn[339]),
.io_parallelIn_340(dataIn[340]),
.io_parallelIn_341(dataIn[341]),
.io_parallelIn_342(dataIn[342]),
.io_parallelIn_343(dataIn[343]),
.io_parallelIn_344(dataIn[344]),
.io_parallelIn_345(dataIn[345]),
.io_parallelIn_346(dataIn[346]),
.io_parallelIn_347(dataIn[347]),
.io_parallelIn_348(dataIn[348]),
.io_parallelIn_349(dataIn[349]),
.io_parallelIn_350(dataIn[350]),
.io_parallelIn_351(dataIn[351]),
.io_parallelIn_352(dataIn[352]),
.io_parallelIn_353(dataIn[353]),
.io_parallelIn_354(dataIn[354]),
.io_parallelIn_355(dataIn[355]),
.io_parallelIn_356(dataIn[356]),
.io_parallelIn_357(dataIn[357]),
.io_parallelIn_358(dataIn[358]),
.io_parallelIn_359(dataIn[359]),
.io_parallelIn_360(dataIn[360]),
.io_parallelIn_361(dataIn[361]),
.io_parallelIn_362(dataIn[362]),
.io_parallelIn_363(dataIn[363]),
.io_parallelIn_364(dataIn[364]),
.io_parallelIn_365(dataIn[365]),
.io_parallelIn_366(dataIn[366]),
.io_parallelIn_367(dataIn[367]),
.io_parallelIn_368(dataIn[368]),
.io_parallelIn_369(dataIn[369]),
.io_parallelIn_370(dataIn[370]),
.io_parallelIn_371(dataIn[371]),
.io_parallelIn_372(dataIn[372]),
.io_parallelIn_373(dataIn[373]),
.io_parallelIn_374(dataIn[374]),
.io_parallelIn_375(dataIn[375]),
.io_parallelIn_376(dataIn[376]),
.io_parallelIn_377(dataIn[377]),
.io_parallelIn_378(dataIn[378]),
.io_parallelIn_379(dataIn[379]),
.io_parallelIn_380(dataIn[380]),
.io_parallelIn_381(dataIn[381]),
.io_parallelIn_382(dataIn[382]),
.io_parallelIn_383(dataIn[383]),
.io_parallelIn_384(dataIn[384]),
.io_parallelIn_385(dataIn[385]),
.io_parallelIn_386(dataIn[386]),
.io_parallelIn_387(dataIn[387]),
.io_parallelIn_388(dataIn[388]),
.io_parallelIn_389(dataIn[389]),
.io_parallelIn_390(dataIn[390]),
.io_parallelIn_391(dataIn[391]),
.io_parallelIn_392(dataIn[392]),
.io_parallelIn_393(dataIn[393]),
.io_parallelIn_394(dataIn[394]),
.io_parallelIn_395(dataIn[395]),
.io_parallelIn_396(dataIn[396]),
.io_parallelIn_397(dataIn[397]),
.io_parallelIn_398(dataIn[398]),
.io_parallelIn_399(dataIn[399]),
.io_parallelIn_400(dataIn[400]),
.io_parallelIn_401(dataIn[401]),
.io_parallelIn_402(dataIn[402]),
.io_parallelIn_403(dataIn[403]),
.io_parallelIn_404(dataIn[404]),
.io_parallelIn_405(dataIn[405]),
.io_parallelIn_406(dataIn[406]),
.io_parallelIn_407(dataIn[407]),
.io_parallelIn_408(dataIn[408]),
.io_parallelIn_409(dataIn[409]),
.io_parallelIn_410(dataIn[410]),
.io_parallelIn_411(dataIn[411]),
.io_parallelIn_412(dataIn[412]),
.io_parallelIn_413(dataIn[413]),
.io_parallelIn_414(dataIn[414]),
.io_parallelIn_415(dataIn[415]),
.io_parallelIn_416(dataIn[416]),
.io_parallelIn_417(dataIn[417]),
.io_parallelIn_418(dataIn[418]),
.io_parallelIn_419(dataIn[419]),
.io_parallelIn_420(dataIn[420]),
.io_parallelIn_421(dataIn[421]),
.io_parallelIn_422(dataIn[422]),
.io_parallelIn_423(dataIn[423]),
.io_parallelIn_424(dataIn[424]),
.io_parallelIn_425(dataIn[425]),
.io_parallelIn_426(dataIn[426]),
.io_parallelIn_427(dataIn[427]),
.io_parallelIn_428(dataIn[428]),
.io_parallelIn_429(dataIn[429]),
.io_parallelIn_430(dataIn[430]),
.io_parallelIn_431(dataIn[431]),
.io_parallelIn_432(dataIn[432]),
.io_parallelIn_433(dataIn[433]),
.io_parallelIn_434(dataIn[434]),
.io_parallelIn_435(dataIn[435]),
.io_parallelIn_436(dataIn[436]),
.io_parallelIn_437(dataIn[437]),
.io_parallelIn_438(dataIn[438]),
.io_parallelIn_439(dataIn[439]),
.io_parallelIn_440(dataIn[440]),
.io_parallelIn_441(dataIn[441]),
.io_parallelIn_442(dataIn[442]),
.io_parallelIn_443(dataIn[443]),
.io_parallelIn_444(dataIn[444]),
.io_parallelIn_445(dataIn[445]),
.io_parallelIn_446(dataIn[446]),
.io_parallelIn_447(dataIn[447]),
.io_parallelIn_448(dataIn[448]),
.io_parallelIn_449(dataIn[449]),
.io_parallelIn_450(dataIn[450]),
.io_parallelIn_451(dataIn[451]),
.io_parallelIn_452(dataIn[452]),
.io_parallelIn_453(dataIn[453]),
.io_parallelIn_454(dataIn[454]),
.io_parallelIn_455(dataIn[455]),
.io_parallelIn_456(dataIn[456]),
.io_parallelIn_457(dataIn[457]),
.io_parallelIn_458(dataIn[458]),
.io_parallelIn_459(dataIn[459]),
.io_parallelIn_460(dataIn[460]),
.io_parallelIn_461(dataIn[461]),
.io_parallelIn_462(dataIn[462]),
.io_parallelIn_463(dataIn[463]),
.io_parallelIn_464(dataIn[464]),
.io_parallelIn_465(dataIn[465]),
.io_parallelIn_466(dataIn[466]),
.io_parallelIn_467(dataIn[467]),
.io_parallelIn_468(dataIn[468]),
.io_parallelIn_469(dataIn[469]),
.io_parallelIn_470(dataIn[470]),
.io_parallelIn_471(dataIn[471]),
.io_parallelIn_472(dataIn[472]),
.io_parallelIn_473(dataIn[473]),
.io_parallelIn_474(dataIn[474]),
.io_parallelIn_475(dataIn[475]),
.io_parallelIn_476(dataIn[476]),
.io_parallelIn_477(dataIn[477]),
.io_parallelIn_478(dataIn[478]),
.io_parallelIn_479(dataIn[479]),
.io_parallelIn_480(dataIn[480]),
.io_parallelIn_481(dataIn[481]),
.io_parallelIn_482(dataIn[482]),
.io_parallelIn_483(dataIn[483]),
.io_parallelIn_484(dataIn[484]),
.io_parallelIn_485(dataIn[485]),
.io_parallelIn_486(dataIn[486]),
.io_parallelIn_487(dataIn[487]),
.io_parallelIn_488(dataIn[488]),
.io_parallelIn_489(dataIn[489]),
.io_parallelIn_490(dataIn[490]),
.io_parallelIn_491(dataIn[491]),
.io_parallelIn_492(dataIn[492]),
.io_parallelIn_493(dataIn[493]),
.io_parallelIn_494(dataIn[494]),
.io_parallelIn_495(dataIn[495]),
.io_parallelIn_496(dataIn[496]),
.io_parallelIn_497(dataIn[497]),
.io_parallelIn_498(dataIn[498]),
.io_parallelIn_499(dataIn[499]),
.io_parallelIn_500(dataIn[500]),
.io_parallelIn_501(dataIn[501]),
.io_parallelIn_502(dataIn[502]),
.io_parallelIn_503(dataIn[503]),
.io_parallelIn_504(dataIn[504]),
.io_parallelIn_505(dataIn[505]),
.io_parallelIn_506(dataIn[506]),
.io_parallelIn_507(dataIn[507]),
.io_parallelIn_508(dataIn[508]),
.io_parallelIn_509(dataIn[509]),
.io_parallelIn_510(dataIn[510]),
.io_parallelIn_511(dataIn[511]),
.io_parallelIn_512(dataIn[512]),
.io_parallelIn_513(dataIn[513]),
.io_parallelIn_514(dataIn[514]),
.io_parallelIn_515(dataIn[515]),
.io_parallelIn_516(dataIn[516]),
.io_parallelIn_517(dataIn[517]),
.io_parallelIn_518(dataIn[518]),
.io_parallelIn_519(dataIn[519]),
.io_parallelIn_520(dataIn[520]),
.io_parallelIn_521(dataIn[521]),
.io_parallelIn_522(dataIn[522]),
.io_parallelIn_523(dataIn[523]),
.io_parallelIn_524(dataIn[524]),
.io_parallelIn_525(dataIn[525]),
.io_parallelIn_526(dataIn[526]),
.io_parallelIn_527(dataIn[527]),
.io_parallelIn_528(dataIn[528]),
.io_parallelIn_529(dataIn[529]),
.io_parallelIn_530(dataIn[530]),
.io_parallelIn_531(dataIn[531]),
.io_parallelIn_532(dataIn[532]),
.io_parallelIn_533(dataIn[533]),
.io_parallelIn_534(dataIn[534]),
.io_parallelIn_535(dataIn[535]),
.io_parallelIn_536(dataIn[536]),
.io_parallelIn_537(dataIn[537]),
.io_parallelIn_538(dataIn[538]),
.io_parallelIn_539(dataIn[539]),
.io_parallelIn_540(dataIn[540]),
.io_parallelIn_541(dataIn[541]),
.io_parallelIn_542(dataIn[542]),
.io_parallelIn_543(dataIn[543]),
.io_parallelIn_544(dataIn[544]),
.io_parallelIn_545(dataIn[545]),
.io_parallelIn_546(dataIn[546]),
.io_parallelIn_547(dataIn[547]),
.io_parallelIn_548(dataIn[548]),
.io_parallelIn_549(dataIn[549]),
.io_parallelIn_550(dataIn[550]),
.io_parallelIn_551(dataIn[551]),
.io_parallelIn_552(dataIn[552]),
.io_parallelIn_553(dataIn[553]),
.io_parallelIn_554(dataIn[554]),
.io_parallelIn_555(dataIn[555]),
.io_parallelIn_556(dataIn[556]),
.io_parallelIn_557(dataIn[557]),
.io_parallelIn_558(dataIn[558]),
.io_parallelIn_559(dataIn[559]),
.io_parallelIn_560(dataIn[560]),
.io_parallelIn_561(dataIn[561]),
.io_parallelIn_562(dataIn[562]),
.io_parallelIn_563(dataIn[563]),
.io_parallelIn_564(dataIn[564]),
.io_parallelIn_565(dataIn[565]),
.io_parallelIn_566(dataIn[566]),
.io_parallelIn_567(dataIn[567]),
.io_parallelIn_568(dataIn[568]),
.io_parallelIn_569(dataIn[569]),
.io_parallelIn_570(dataIn[570]),
.io_parallelIn_571(dataIn[571]),
.io_parallelIn_572(dataIn[572]),
.io_parallelIn_573(dataIn[573]),
.io_parallelIn_574(dataIn[574]),
.io_parallelIn_575(dataIn[575]),
.io_parallelIn_576(dataIn[576]),
.io_parallelIn_577(dataIn[577]),
.io_parallelIn_578(dataIn[578]),
.io_parallelIn_579(dataIn[579]),
.io_parallelIn_580(dataIn[580]),
.io_parallelIn_581(dataIn[581]),
.io_parallelIn_582(dataIn[582]),
.io_parallelIn_583(dataIn[583]),
.io_parallelIn_584(dataIn[584]),
.io_parallelIn_585(dataIn[585]),
.io_parallelIn_586(dataIn[586]),
.io_parallelIn_587(dataIn[587]),
.io_parallelIn_588(dataIn[588]),
.io_parallelIn_589(dataIn[589]),
.io_parallelIn_590(dataIn[590]),
.io_parallelIn_591(dataIn[591]),
.io_parallelIn_592(dataIn[592]),
.io_parallelIn_593(dataIn[593]),
.io_parallelIn_594(dataIn[594]),
.io_parallelIn_595(dataIn[595]),
.io_parallelIn_596(dataIn[596]),
.io_parallelIn_597(dataIn[597]),
.io_parallelIn_598(dataIn[598]),
.io_parallelIn_599(dataIn[599]),
.io_parallelIn_600(dataIn[600]),
.io_parallelIn_601(dataIn[601]),
.io_parallelIn_602(dataIn[602]),
.io_parallelIn_603(dataIn[603]),
.io_parallelIn_604(dataIn[604]),
.io_parallelIn_605(dataIn[605]),
.io_parallelIn_606(dataIn[606]),
.io_parallelIn_607(dataIn[607]),
.io_parallelIn_608(dataIn[608]),
.io_parallelIn_609(dataIn[609]),
.io_parallelIn_610(dataIn[610]),
.io_parallelIn_611(dataIn[611]),
.io_parallelIn_612(dataIn[612]),
.io_parallelIn_613(dataIn[613]),
.io_parallelIn_614(dataIn[614]),
.io_parallelIn_615(dataIn[615]),
.io_parallelIn_616(dataIn[616]),
.io_parallelIn_617(dataIn[617]),
.io_parallelIn_618(dataIn[618]),
.io_parallelIn_619(dataIn[619]),
.io_parallelIn_620(dataIn[620]),
.io_parallelIn_621(dataIn[621]),
.io_parallelIn_622(dataIn[622]),
.io_parallelIn_623(dataIn[623]),
.io_parallelIn_624(dataIn[624]),
.io_parallelIn_625(dataIn[625]),
.io_parallelIn_626(dataIn[626]),
.io_parallelIn_627(dataIn[627]),
.io_parallelIn_628(dataIn[628]),
.io_parallelIn_629(dataIn[629]),
.io_parallelIn_630(dataIn[630]),
.io_parallelIn_631(dataIn[631]),
.io_parallelIn_632(dataIn[632]),
.io_parallelIn_633(dataIn[633]),
.io_parallelIn_634(dataIn[634]),
.io_parallelIn_635(dataIn[635]),
.io_parallelIn_636(dataIn[636]),
.io_parallelIn_637(dataIn[637]),
.io_parallelIn_638(dataIn[638]),
.io_parallelIn_639(dataIn[639]),
.io_parallelIn_640(dataIn[640]),
.io_parallelIn_641(dataIn[641]),
.io_parallelIn_642(dataIn[642]),
.io_parallelIn_643(dataIn[643]),
.io_parallelIn_644(dataIn[644]),
.io_parallelIn_645(dataIn[645]),
.io_parallelIn_646(dataIn[646]),
.io_parallelIn_647(dataIn[647]),
.io_parallelIn_648(dataIn[648]),
.io_parallelIn_649(dataIn[649]),
.io_parallelIn_650(dataIn[650]),
.io_parallelIn_651(dataIn[651]),
.io_parallelIn_652(dataIn[652]),
.io_parallelIn_653(dataIn[653]),
.io_parallelIn_654(dataIn[654]),
.io_parallelIn_655(dataIn[655]),
.io_parallelIn_656(dataIn[656]),
.io_parallelIn_657(dataIn[657]),
.io_parallelIn_658(dataIn[658]),
.io_parallelIn_659(dataIn[659]),
.io_parallelIn_660(dataIn[660]),
.io_parallelIn_661(dataIn[661]),
.io_parallelIn_662(dataIn[662]),
.io_parallelIn_663(dataIn[663]),
.io_parallelIn_664(dataIn[664]),
.io_parallelIn_665(dataIn[665]),
.io_parallelIn_666(dataIn[666]),
.io_parallelIn_667(dataIn[667]),
.io_parallelIn_668(dataIn[668]),
.io_parallelIn_669(dataIn[669]),
.io_parallelIn_670(dataIn[670]),
.io_parallelIn_671(dataIn[671]),
.io_parallelIn_672(dataIn[672]),
.io_parallelIn_673(dataIn[673]),
.io_parallelIn_674(dataIn[674]),
.io_parallelIn_675(dataIn[675]),
.io_parallelIn_676(dataIn[676]),
.io_parallelIn_677(dataIn[677]),
.io_parallelIn_678(dataIn[678]),
.io_parallelIn_679(dataIn[679]),
.io_parallelIn_680(dataIn[680]),
.io_parallelIn_681(dataIn[681]),
.io_parallelIn_682(dataIn[682]),
.io_parallelIn_683(dataIn[683]),
.io_parallelIn_684(dataIn[684]),
.io_parallelIn_685(dataIn[685]),
.io_parallelIn_686(dataIn[686]),
.io_parallelIn_687(dataIn[687]),
.io_parallelIn_688(dataIn[688]),
.io_parallelIn_689(dataIn[689]),
.io_parallelIn_690(dataIn[690]),
.io_parallelIn_691(dataIn[691]),
.io_parallelIn_692(dataIn[692]),
.io_parallelIn_693(dataIn[693]),
.io_parallelIn_694(dataIn[694]),
.io_parallelIn_695(dataIn[695]),
.io_parallelIn_696(dataIn[696]),
.io_parallelIn_697(dataIn[697]),
.io_parallelIn_698(dataIn[698]),
.io_parallelIn_699(dataIn[699]),
.io_parallelIn_700(dataIn[700]),
.io_parallelIn_701(dataIn[701]),
.io_parallelIn_702(dataIn[702]),
.io_parallelIn_703(dataIn[703]),
.io_parallelIn_704(dataIn[704]),
.io_parallelIn_705(dataIn[705]),
.io_parallelIn_706(dataIn[706]),
.io_parallelIn_707(dataIn[707]),
.io_parallelIn_708(dataIn[708]),
.io_parallelIn_709(dataIn[709]),
.io_parallelIn_710(dataIn[710]),
.io_parallelIn_711(dataIn[711]),
.io_parallelIn_712(dataIn[712]),
.io_parallelIn_713(dataIn[713]),
.io_parallelIn_714(dataIn[714]),
.io_parallelIn_715(dataIn[715]),
.io_parallelIn_716(dataIn[716]),
.io_parallelIn_717(dataIn[717]),
.io_parallelIn_718(dataIn[718]),
.io_parallelIn_719(dataIn[719]),
.io_parallelIn_720(dataIn[720]),
.io_parallelIn_721(dataIn[721]),
.io_parallelIn_722(dataIn[722]),
.io_parallelIn_723(dataIn[723]),
.io_parallelIn_724(dataIn[724]),
.io_parallelIn_725(dataIn[725]),
.io_parallelIn_726(dataIn[726]),
.io_parallelIn_727(dataIn[727]),
.io_parallelIn_728(dataIn[728]),
.io_parallelIn_729(dataIn[729]),
.io_parallelIn_730(dataIn[730]),
.io_parallelIn_731(dataIn[731]),
.io_parallelIn_732(dataIn[732]),
.io_parallelIn_733(dataIn[733]),
.io_parallelIn_734(dataIn[734]),
.io_parallelIn_735(dataIn[735]),
.io_parallelIn_736(dataIn[736]),
.io_parallelIn_737(dataIn[737]),
.io_parallelIn_738(dataIn[738]),
.io_parallelIn_739(dataIn[739]),
.io_parallelIn_740(dataIn[740]),
.io_parallelIn_741(dataIn[741]),
.io_parallelIn_742(dataIn[742]),
.io_parallelIn_743(dataIn[743]),
.io_parallelIn_744(dataIn[744]),
.io_parallelIn_745(dataIn[745]),
.io_parallelIn_746(dataIn[746]),
.io_parallelIn_747(dataIn[747]),
.io_parallelIn_748(dataIn[748]),
.io_parallelIn_749(dataIn[749]),
.io_parallelIn_750(dataIn[750]),
.io_parallelIn_751(dataIn[751]),
.io_parallelIn_752(dataIn[752]),
.io_parallelIn_753(dataIn[753]),
.io_parallelIn_754(dataIn[754]),
.io_parallelIn_755(dataIn[755]),
.io_parallelIn_756(dataIn[756]),
.io_parallelIn_757(dataIn[757]),
.io_parallelIn_758(dataIn[758]),
.io_parallelIn_759(dataIn[759]),
.io_parallelIn_760(dataIn[760]),
.io_parallelIn_761(dataIn[761]),
.io_parallelIn_762(dataIn[762]),
.io_parallelIn_763(dataIn[763]),
.io_parallelIn_764(dataIn[764]),
.io_parallelIn_765(dataIn[765]),
.io_parallelIn_766(dataIn[766]),
.io_parallelIn_767(dataIn[767]),
.io_parallelIn_768(dataIn[768]),
.io_parallelIn_769(dataIn[769]),
.io_parallelIn_770(dataIn[770]),
.io_parallelIn_771(dataIn[771]),
.io_parallelIn_772(dataIn[772]),
.io_parallelIn_773(dataIn[773]),
.io_parallelIn_774(dataIn[774]),
.io_parallelIn_775(dataIn[775]),
.io_parallelIn_776(dataIn[776]),
.io_parallelIn_777(dataIn[777]),
.io_parallelIn_778(dataIn[778]),
.io_parallelIn_779(dataIn[779]),
.io_parallelIn_780(dataIn[780]),
.io_parallelIn_781(dataIn[781]),
.io_parallelIn_782(dataIn[782]),
.io_parallelIn_783(dataIn[783]),
.io_parallelIn_784(dataIn[784]),
.io_parallelIn_785(dataIn[785]),
.io_parallelIn_786(dataIn[786]),
.io_parallelIn_787(dataIn[787]),
.io_parallelIn_788(dataIn[788]),
.io_parallelIn_789(dataIn[789]),
.io_parallelIn_790(dataIn[790]),
.io_parallelIn_791(dataIn[791]),
.io_parallelIn_792(dataIn[792]),
.io_parallelIn_793(dataIn[793]),
.io_parallelIn_794(dataIn[794]),
.io_parallelIn_795(dataIn[795]),
.io_parallelIn_796(dataIn[796]),
.io_parallelIn_797(dataIn[797]),
.io_parallelIn_798(dataIn[798]),
.io_parallelIn_799(dataIn[799]),
.io_parallelIn_800(dataIn[800]),
.io_parallelIn_801(dataIn[801]),
.io_parallelIn_802(dataIn[802]),
.io_parallelIn_803(dataIn[803]),
.io_parallelIn_804(dataIn[804]),
.io_parallelIn_805(dataIn[805]),
.io_parallelIn_806(dataIn[806]),
.io_parallelIn_807(dataIn[807]),
.io_parallelIn_808(dataIn[808]),
.io_parallelIn_809(dataIn[809]),
.io_parallelIn_810(dataIn[810]),
.io_parallelIn_811(dataIn[811]),
.io_parallelIn_812(dataIn[812]),
.io_parallelIn_813(dataIn[813]),
.io_parallelIn_814(dataIn[814]),
.io_parallelIn_815(dataIn[815]),
.io_parallelIn_816(dataIn[816]),
.io_parallelIn_817(dataIn[817]),
.io_parallelIn_818(dataIn[818]),
.io_parallelIn_819(dataIn[819]),
.io_parallelIn_820(dataIn[820]),
.io_parallelIn_821(dataIn[821]),
.io_parallelIn_822(dataIn[822]),
.io_parallelIn_823(dataIn[823]),
.io_parallelIn_824(dataIn[824]),
.io_parallelIn_825(dataIn[825]),
.io_parallelIn_826(dataIn[826]),
.io_parallelIn_827(dataIn[827]),
.io_parallelIn_828(dataIn[828]),
.io_parallelIn_829(dataIn[829]),
.io_parallelIn_830(dataIn[830]),
.io_parallelIn_831(dataIn[831]),
.io_parallelIn_832(dataIn[832]),
.io_parallelIn_833(dataIn[833]),
.io_parallelIn_834(dataIn[834]),
.io_parallelIn_835(dataIn[835]),
.io_parallelIn_836(dataIn[836]),
.io_parallelIn_837(dataIn[837]),
.io_parallelIn_838(dataIn[838]),
.io_parallelIn_839(dataIn[839]),
.io_parallelIn_840(dataIn[840]),
.io_parallelIn_841(dataIn[841]),
.io_parallelIn_842(dataIn[842]),
.io_parallelIn_843(dataIn[843]),
.io_parallelIn_844(dataIn[844]),
.io_parallelIn_845(dataIn[845]),
.io_parallelIn_846(dataIn[846]),
.io_parallelIn_847(dataIn[847]),
.io_parallelIn_848(dataIn[848]),
.io_parallelIn_849(dataIn[849]),
.io_parallelIn_850(dataIn[850]),
.io_parallelIn_851(dataIn[851]),
.io_parallelIn_852(dataIn[852]),
.io_parallelIn_853(dataIn[853]),
.io_parallelIn_854(dataIn[854]),
.io_parallelIn_855(dataIn[855]),
.io_parallelIn_856(dataIn[856]),
.io_parallelIn_857(dataIn[857]),
.io_parallelIn_858(dataIn[858]),
.io_parallelIn_859(dataIn[859]),
.io_parallelIn_860(dataIn[860]),
.io_parallelIn_861(dataIn[861]),
.io_parallelIn_862(dataIn[862]),
.io_parallelIn_863(dataIn[863]),
.io_parallelIn_864(dataIn[864]),
.io_parallelIn_865(dataIn[865]),
.io_parallelIn_866(dataIn[866]),
.io_parallelIn_867(dataIn[867]),
.io_parallelIn_868(dataIn[868]),
.io_parallelIn_869(dataIn[869]),
.io_parallelIn_870(dataIn[870]),
.io_parallelIn_871(dataIn[871]),
.io_parallelIn_872(dataIn[872]),
.io_parallelIn_873(dataIn[873]),
.io_parallelIn_874(dataIn[874]),
.io_parallelIn_875(dataIn[875]),
.io_parallelIn_876(dataIn[876]),
.io_parallelIn_877(dataIn[877]),
.io_parallelIn_878(dataIn[878]),
.io_parallelIn_879(dataIn[879]),
.io_parallelIn_880(dataIn[880]),
.io_parallelIn_881(dataIn[881]),
.io_parallelIn_882(dataIn[882]),
.io_parallelIn_883(dataIn[883]),
.io_parallelIn_884(dataIn[884]),
.io_parallelIn_885(dataIn[885]),
.io_parallelIn_886(dataIn[886]),
.io_parallelIn_887(dataIn[887]),
.io_parallelIn_888(dataIn[888]),
.io_parallelIn_889(dataIn[889]),
.io_parallelIn_890(dataIn[890]),
.io_parallelIn_891(dataIn[891]),
.io_parallelIn_892(dataIn[892]),
.io_parallelIn_893(dataIn[893]),
.io_parallelIn_894(dataIn[894]),
.io_parallelIn_895(dataIn[895]),
.io_parallelIn_896(dataIn[896]),
.io_parallelIn_897(dataIn[897]),
.io_parallelIn_898(dataIn[898]),
.io_parallelIn_899(dataIn[899]),
.io_parallelIn_900(dataIn[900]),
.io_parallelIn_901(dataIn[901]),
.io_parallelIn_902(dataIn[902]),
.io_parallelIn_903(dataIn[903]),
.io_parallelIn_904(dataIn[904]),
.io_parallelIn_905(dataIn[905]),
.io_parallelIn_906(dataIn[906]),
.io_parallelIn_907(dataIn[907]),
.io_parallelIn_908(dataIn[908]),
.io_parallelIn_909(dataIn[909]),
.io_parallelIn_910(dataIn[910]),
.io_parallelIn_911(dataIn[911]),
.io_parallelIn_912(dataIn[912]),
.io_parallelIn_913(dataIn[913]),
.io_parallelIn_914(dataIn[914]),
.io_parallelIn_915(dataIn[915]),
.io_parallelIn_916(dataIn[916]),
.io_parallelIn_917(dataIn[917]),
.io_parallelIn_918(dataIn[918]),
.io_parallelIn_919(dataIn[919]),
.io_parallelIn_920(dataIn[920]),
.io_parallelIn_921(dataIn[921]),
.io_parallelIn_922(dataIn[922]),
.io_parallelIn_923(dataIn[923]),
.io_parallelIn_924(dataIn[924]),
.io_parallelIn_925(dataIn[925]),
.io_parallelIn_926(dataIn[926]),
.io_parallelIn_927(dataIn[927]),
.io_parallelIn_928(dataIn[928]),
.io_parallelIn_929(dataIn[929]),
.io_parallelIn_930(dataIn[930]),
.io_parallelIn_931(dataIn[931]),
.io_parallelIn_932(dataIn[932]),
.io_parallelIn_933(dataIn[933]),
.io_parallelIn_934(dataIn[934]),
.io_parallelIn_935(dataIn[935]),
.io_parallelIn_936(dataIn[936]),
.io_parallelIn_937(dataIn[937]),
.io_parallelIn_938(dataIn[938]),
.io_parallelIn_939(dataIn[939]),
.io_parallelIn_940(dataIn[940]),
.io_parallelIn_941(dataIn[941]),
.io_parallelIn_942(dataIn[942]),
.io_parallelIn_943(dataIn[943]),
.io_parallelIn_944(dataIn[944]),
.io_parallelIn_945(dataIn[945]),
.io_parallelIn_946(dataIn[946]),
.io_parallelIn_947(dataIn[947]),
.io_parallelIn_948(dataIn[948]),
.io_parallelIn_949(dataIn[949]),
.io_parallelIn_950(dataIn[950]),
.io_parallelIn_951(dataIn[951]),
.io_parallelIn_952(dataIn[952]),
.io_parallelIn_953(dataIn[953]),
.io_parallelIn_954(dataIn[954]),
.io_parallelIn_955(dataIn[955]),
.io_parallelIn_956(dataIn[956]),
.io_parallelIn_957(dataIn[957]),
.io_parallelIn_958(dataIn[958]),
.io_parallelIn_959(dataIn[959]),
.io_parallelIn_960(dataIn[960]),
.io_parallelIn_961(dataIn[961]),
.io_parallelIn_962(dataIn[962]),
.io_parallelIn_963(dataIn[963]),
.io_parallelIn_964(dataIn[964]),
.io_parallelIn_965(dataIn[965]),
.io_parallelIn_966(dataIn[966]),
.io_parallelIn_967(dataIn[967]),
.io_parallelIn_968(dataIn[968]),
.io_parallelIn_969(dataIn[969]),
.io_parallelIn_970(dataIn[970]),
.io_parallelIn_971(dataIn[971]),
.io_parallelIn_972(dataIn[972]),
.io_parallelIn_973(dataIn[973]),
.io_parallelIn_974(dataIn[974]),
.io_parallelIn_975(dataIn[975]),
.io_parallelIn_976(dataIn[976]),
.io_parallelIn_977(dataIn[977]),
.io_parallelIn_978(dataIn[978]),
.io_parallelIn_979(dataIn[979]),
.io_parallelIn_980(dataIn[980]),
.io_parallelIn_981(dataIn[981]),
.io_parallelIn_982(dataIn[982]),
.io_parallelIn_983(dataIn[983]),
.io_parallelIn_984(dataIn[984]),
.io_parallelIn_985(dataIn[985]),
.io_parallelIn_986(dataIn[986]),
.io_parallelIn_987(dataIn[987]),
.io_parallelIn_988(dataIn[988]),
.io_parallelIn_989(dataIn[989]),
.io_parallelIn_990(dataIn[990]),
.io_parallelIn_991(dataIn[991]),
.io_parallelIn_992(dataIn[992]),
.io_parallelIn_993(dataIn[993]),
.io_parallelIn_994(dataIn[994]),
.io_parallelIn_995(dataIn[995]),
.io_parallelIn_996(dataIn[996]),
.io_parallelIn_997(dataIn[997]),
.io_parallelIn_998(dataIn[998]),
.io_parallelIn_999(dataIn[999]),
.io_parallelIn_1000(dataIn[1000]),
.io_parallelIn_1001(dataIn[1001]),
.io_parallelIn_1002(dataIn[1002]),
.io_parallelIn_1003(dataIn[1003]),
.io_parallelIn_1004(dataIn[1004]),
.io_parallelIn_1005(dataIn[1005]),
.io_parallelIn_1006(dataIn[1006]),
.io_parallelIn_1007(dataIn[1007]),
.io_parallelIn_1008(dataIn[1008]),
.io_parallelIn_1009(dataIn[1009]),
.io_parallelIn_1010(dataIn[1010]),
.io_parallelIn_1011(dataIn[1011]),
.io_parallelIn_1012(dataIn[1012]),
.io_parallelIn_1013(dataIn[1013]),
.io_parallelIn_1014(dataIn[1014]),
.io_parallelIn_1015(dataIn[1015]),
.io_parallelIn_1016(dataIn[1016]),
.io_parallelIn_1017(dataIn[1017]),
.io_parallelIn_1018(dataIn[1018]),
.io_parallelIn_1019(dataIn[1019]),
.io_parallelIn_1020(dataIn[1020]),
.io_parallelIn_1021(dataIn[1021]),
.io_parallelIn_1022(dataIn[1022]),
.io_parallelIn_1023(dataIn[1023]),
.io_parallelIn_1024(dataIn[1024]),
.io_parallelIn_1025(dataIn[1025]),
.io_parallelIn_1026(dataIn[1026]),
.io_parallelIn_1027(dataIn[1027]),
.io_parallelIn_1028(dataIn[1028]),
.io_parallelIn_1029(dataIn[1029]),
.io_parallelIn_1030(dataIn[1030]),
.io_parallelIn_1031(dataIn[1031]),
.io_parallelIn_1032(dataIn[1032]),
.io_parallelIn_1033(dataIn[1033]),
.io_parallelIn_1034(dataIn[1034]),
.io_parallelIn_1035(dataIn[1035]),
.io_parallelIn_1036(dataIn[1036]),
.io_parallelIn_1037(dataIn[1037]),
.io_parallelIn_1038(dataIn[1038]),
.io_parallelIn_1039(dataIn[1039]),
.io_parallelIn_1040(dataIn[1040]),
.io_parallelIn_1041(dataIn[1041]),
.io_parallelIn_1042(dataIn[1042]),
.io_parallelIn_1043(dataIn[1043]),
.io_parallelIn_1044(dataIn[1044]),
.io_parallelIn_1045(dataIn[1045]),
.io_parallelIn_1046(dataIn[1046]),
.io_parallelIn_1047(dataIn[1047]),
.io_parallelIn_1048(dataIn[1048]),
.io_parallelIn_1049(dataIn[1049]),
.io_parallelIn_1050(dataIn[1050]),
.io_parallelIn_1051(dataIn[1051]),
.io_parallelIn_1052(dataIn[1052]),
.io_parallelIn_1053(dataIn[1053]),
.io_parallelIn_1054(dataIn[1054]),
.io_parallelIn_1055(dataIn[1055]),
.io_parallelIn_1056(dataIn[1056]),
.io_parallelIn_1057(dataIn[1057]),
.io_parallelIn_1058(dataIn[1058]),
.io_parallelIn_1059(dataIn[1059]),
.io_parallelIn_1060(dataIn[1060]),
.io_parallelIn_1061(dataIn[1061]),
.io_parallelIn_1062(dataIn[1062]),
.io_parallelIn_1063(dataIn[1063]),
.io_parallelIn_1064(dataIn[1064]),
.io_parallelIn_1065(dataIn[1065]),
.io_parallelIn_1066(dataIn[1066]),
.io_parallelIn_1067(dataIn[1067]),
.io_parallelIn_1068(dataIn[1068]),
.io_parallelIn_1069(dataIn[1069]),
.io_parallelIn_1070(dataIn[1070]),
.io_parallelIn_1071(dataIn[1071]),
.io_parallelIn_1072(dataIn[1072]),
.io_parallelIn_1073(dataIn[1073]),
.io_parallelIn_1074(dataIn[1074]),
.io_parallelIn_1075(dataIn[1075]),
.io_parallelIn_1076(dataIn[1076]),
.io_parallelIn_1077(dataIn[1077]),
.io_parallelIn_1078(dataIn[1078]),
.io_parallelIn_1079(dataIn[1079]),
.io_parallelIn_1080(dataIn[1080]),
.io_parallelIn_1081(dataIn[1081]),
.io_parallelIn_1082(dataIn[1082]),
.io_parallelIn_1083(dataIn[1083]),
.io_parallelIn_1084(dataIn[1084]),
.io_parallelIn_1085(dataIn[1085]),
.io_parallelIn_1086(dataIn[1086]),
.io_parallelIn_1087(dataIn[1087]),
.io_parallelIn_1088(dataIn[1088]),
.io_parallelIn_1089(dataIn[1089]),
.io_parallelIn_1090(dataIn[1090]),
.io_parallelIn_1091(dataIn[1091]),
.io_parallelIn_1092(dataIn[1092]),
.io_parallelIn_1093(dataIn[1093]),
.io_parallelIn_1094(dataIn[1094]),
.io_parallelIn_1095(dataIn[1095]),
.io_parallelIn_1096(dataIn[1096]),
.io_parallelIn_1097(dataIn[1097]),
.io_parallelIn_1098(dataIn[1098]),
.io_parallelIn_1099(dataIn[1099]),
.io_parallelIn_1100(dataIn[1100]),
.io_parallelIn_1101(dataIn[1101]),
.io_parallelIn_1102(dataIn[1102]),
.io_parallelIn_1103(dataIn[1103]),
.io_parallelIn_1104(dataIn[1104]),
.io_parallelIn_1105(dataIn[1105]),
.io_parallelIn_1106(dataIn[1106]),
.io_parallelIn_1107(dataIn[1107]),
.io_parallelIn_1108(dataIn[1108]),
.io_parallelIn_1109(dataIn[1109]),
.io_parallelIn_1110(dataIn[1110]),
.io_parallelIn_1111(dataIn[1111]),
.io_parallelIn_1112(dataIn[1112]),
.io_parallelIn_1113(dataIn[1113]),
.io_parallelIn_1114(dataIn[1114]),
.io_parallelIn_1115(dataIn[1115]),
.io_parallelIn_1116(dataIn[1116]),
.io_parallelIn_1117(dataIn[1117]),
.io_parallelIn_1118(dataIn[1118]),
.io_parallelIn_1119(dataIn[1119]),
.io_parallelIn_1120(dataIn[1120]),
.io_parallelIn_1121(dataIn[1121]),
.io_parallelIn_1122(dataIn[1122]),
.io_parallelIn_1123(dataIn[1123]),
.io_parallelIn_1124(dataIn[1124]),
.io_parallelIn_1125(dataIn[1125]),
.io_parallelIn_1126(dataIn[1126]),
.io_parallelIn_1127(dataIn[1127]),
.io_parallelIn_1128(dataIn[1128]),
.io_parallelIn_1129(dataIn[1129]),
.io_parallelIn_1130(dataIn[1130]),
.io_parallelIn_1131(dataIn[1131]),
.io_parallelIn_1132(dataIn[1132]),
.io_parallelIn_1133(dataIn[1133]),
.io_parallelIn_1134(dataIn[1134]),
.io_parallelIn_1135(dataIn[1135]),
.io_parallelIn_1136(dataIn[1136]),
.io_parallelIn_1137(dataIn[1137]),
.io_parallelIn_1138(dataIn[1138]),
.io_parallelIn_1139(dataIn[1139]),
.io_parallelIn_1140(dataIn[1140]),
.io_parallelIn_1141(dataIn[1141]),
.io_parallelIn_1142(dataIn[1142]),
.io_parallelIn_1143(dataIn[1143]),
.io_parallelIn_1144(dataIn[1144]),
.io_parallelIn_1145(dataIn[1145]),
.io_parallelIn_1146(dataIn[1146]),
.io_parallelIn_1147(dataIn[1147]),
.io_parallelIn_1148(dataIn[1148]),
.io_parallelIn_1149(dataIn[1149]),
.io_parallelIn_1150(dataIn[1150]),
.io_parallelIn_1151(dataIn[1151]),
.io_parallelIn_1152(dataIn[1152]),
.io_parallelIn_1153(dataIn[1153]),
.io_parallelIn_1154(dataIn[1154]),
.io_parallelIn_1155(dataIn[1155]),
.io_parallelIn_1156(dataIn[1156]),
.io_parallelIn_1157(dataIn[1157]),
.io_parallelIn_1158(dataIn[1158]),
.io_parallelIn_1159(dataIn[1159]),
.io_parallelIn_1160(dataIn[1160]),
.io_parallelIn_1161(dataIn[1161]),
.io_parallelIn_1162(dataIn[1162]),
.io_parallelIn_1163(dataIn[1163]),
.io_parallelIn_1164(dataIn[1164]),
.io_parallelIn_1165(dataIn[1165]),
.io_parallelIn_1166(dataIn[1166]),
.io_parallelIn_1167(dataIn[1167]),
.io_parallelIn_1168(dataIn[1168]),
.io_parallelIn_1169(dataIn[1169]),
.io_parallelIn_1170(dataIn[1170]),
.io_parallelIn_1171(dataIn[1171]),
.io_parallelIn_1172(dataIn[1172]),
.io_parallelIn_1173(dataIn[1173]),
.io_parallelIn_1174(dataIn[1174]),
.io_parallelIn_1175(dataIn[1175]),
.io_parallelIn_1176(dataIn[1176]),
.io_parallelIn_1177(dataIn[1177]),
.io_parallelIn_1178(dataIn[1178]),
.io_parallelIn_1179(dataIn[1179]),
.io_parallelIn_1180(dataIn[1180]),
.io_parallelIn_1181(dataIn[1181]),
.io_parallelIn_1182(dataIn[1182]),
.io_parallelIn_1183(dataIn[1183]),
.io_parallelIn_1184(dataIn[1184]),
.io_parallelIn_1185(dataIn[1185]),
.io_parallelIn_1186(dataIn[1186]),
.io_parallelIn_1187(dataIn[1187]),
.io_parallelIn_1188(dataIn[1188]),
.io_parallelIn_1189(dataIn[1189]),
.io_parallelIn_1190(dataIn[1190]),
.io_parallelIn_1191(dataIn[1191]),
.io_parallelIn_1192(dataIn[1192]),
.io_parallelIn_1193(dataIn[1193]),
.io_parallelIn_1194(dataIn[1194]),
.io_parallelIn_1195(dataIn[1195]),
.io_parallelIn_1196(dataIn[1196]),
.io_parallelIn_1197(dataIn[1197]),
.io_parallelIn_1198(dataIn[1198]),
.io_parallelIn_1199(dataIn[1199]),
.io_parallelIn_1200(dataIn[1200]),
.io_parallelIn_1201(dataIn[1201]),
.io_parallelIn_1202(dataIn[1202]),
.io_parallelIn_1203(dataIn[1203]),
.io_parallelIn_1204(dataIn[1204]),
.io_parallelIn_1205(dataIn[1205]),
.io_parallelIn_1206(dataIn[1206]),
.io_parallelIn_1207(dataIn[1207]),
.io_parallelIn_1208(dataIn[1208]),
.io_parallelIn_1209(dataIn[1209]),
.io_parallelIn_1210(dataIn[1210]),
.io_parallelIn_1211(dataIn[1211]),
.io_parallelIn_1212(dataIn[1212]),
.io_parallelIn_1213(dataIn[1213]),
.io_parallelIn_1214(dataIn[1214]),
.io_parallelIn_1215(dataIn[1215]),
.io_parallelIn_1216(dataIn[1216]),
.io_parallelIn_1217(dataIn[1217]),
.io_parallelIn_1218(dataIn[1218]),
.io_parallelIn_1219(dataIn[1219]),
.io_parallelIn_1220(dataIn[1220]),
.io_parallelIn_1221(dataIn[1221]),
.io_parallelIn_1222(dataIn[1222]),
.io_parallelIn_1223(dataIn[1223]),
.io_parallelIn_1224(dataIn[1224]),
.io_parallelIn_1225(dataIn[1225]),
.io_parallelIn_1226(dataIn[1226]),
.io_parallelIn_1227(dataIn[1227]),
.io_parallelIn_1228(dataIn[1228]),
.io_parallelIn_1229(dataIn[1229]),
.io_parallelIn_1230(dataIn[1230]),
.io_parallelIn_1231(dataIn[1231]),
.io_parallelIn_1232(dataIn[1232]),
.io_parallelIn_1233(dataIn[1233]),
.io_parallelIn_1234(dataIn[1234]),
.io_parallelIn_1235(dataIn[1235]),
.io_parallelIn_1236(dataIn[1236]),
.io_parallelIn_1237(dataIn[1237]),
.io_parallelIn_1238(dataIn[1238]),
.io_parallelIn_1239(dataIn[1239]),
.io_parallelIn_1240(dataIn[1240]),
.io_parallelIn_1241(dataIn[1241]),
.io_parallelIn_1242(dataIn[1242]),
.io_parallelIn_1243(dataIn[1243]),
.io_parallelIn_1244(dataIn[1244]),
.io_parallelIn_1245(dataIn[1245]),
.io_parallelIn_1246(dataIn[1246]),
.io_parallelIn_1247(dataIn[1247]),
.io_parallelIn_1248(dataIn[1248]),
.io_parallelIn_1249(dataIn[1249]),
.io_parallelIn_1250(dataIn[1250]),
.io_parallelIn_1251(dataIn[1251]),
.io_parallelIn_1252(dataIn[1252]),
.io_parallelIn_1253(dataIn[1253]),
.io_parallelIn_1254(dataIn[1254]),
.io_parallelIn_1255(dataIn[1255]),
.io_parallelIn_1256(dataIn[1256]),
.io_parallelIn_1257(dataIn[1257]),
.io_parallelIn_1258(dataIn[1258]),
.io_parallelIn_1259(dataIn[1259]),
.io_parallelIn_1260(dataIn[1260]),
.io_parallelIn_1261(dataIn[1261]),
.io_parallelIn_1262(dataIn[1262]),
.io_parallelIn_1263(dataIn[1263]),
.io_parallelIn_1264(dataIn[1264]),
.io_parallelIn_1265(dataIn[1265]),
.io_parallelIn_1266(dataIn[1266]),
.io_parallelIn_1267(dataIn[1267]),
.io_parallelIn_1268(dataIn[1268]),
.io_parallelIn_1269(dataIn[1269]),
.io_parallelIn_1270(dataIn[1270]),
.io_parallelIn_1271(dataIn[1271]),
.io_parallelIn_1272(dataIn[1272]),
.io_parallelIn_1273(dataIn[1273]),
.io_parallelIn_1274(dataIn[1274]),
.io_parallelIn_1275(dataIn[1275]),
.io_parallelIn_1276(dataIn[1276]),
.io_parallelIn_1277(dataIn[1277]),
.io_parallelIn_1278(dataIn[1278]),
.io_parallelIn_1279(dataIn[1279]),
.io_parallelIn_1280(dataIn[1280]),
.io_parallelIn_1281(dataIn[1281]),
.io_parallelIn_1282(dataIn[1282]),
.io_parallelIn_1283(dataIn[1283]),
.io_parallelIn_1284(dataIn[1284]),
.io_parallelIn_1285(dataIn[1285]),
.io_parallelIn_1286(dataIn[1286]),
.io_parallelIn_1287(dataIn[1287]),
.io_parallelIn_1288(dataIn[1288]),
.io_parallelIn_1289(dataIn[1289]),
.io_parallelIn_1290(dataIn[1290]),
.io_parallelIn_1291(dataIn[1291]),
.io_parallelIn_1292(dataIn[1292]),
.io_parallelIn_1293(dataIn[1293]),
.io_parallelIn_1294(dataIn[1294]),
.io_parallelIn_1295(dataIn[1295]),
.io_parallelIn_1296(dataIn[1296]),
.io_parallelIn_1297(dataIn[1297]),
.io_parallelIn_1298(dataIn[1298]),
.io_parallelIn_1299(dataIn[1299]),
.io_parallelIn_1300(dataIn[1300]),
.io_parallelIn_1301(dataIn[1301]),
.io_parallelIn_1302(dataIn[1302]),
.io_parallelIn_1303(dataIn[1303]),
.io_parallelIn_1304(dataIn[1304]),
.io_parallelIn_1305(dataIn[1305]),
.io_parallelIn_1306(dataIn[1306]),
.io_parallelIn_1307(dataIn[1307]),
.io_parallelIn_1308(dataIn[1308]),
.io_parallelIn_1309(dataIn[1309]),
.io_parallelIn_1310(dataIn[1310]),
.io_parallelIn_1311(dataIn[1311]),
.io_parallelIn_1312(dataIn[1312]),
.io_parallelIn_1313(dataIn[1313]),
.io_parallelIn_1314(dataIn[1314]),
.io_parallelIn_1315(dataIn[1315]),
.io_parallelIn_1316(dataIn[1316]),
.io_parallelIn_1317(dataIn[1317]),
.io_parallelIn_1318(dataIn[1318]),
.io_parallelIn_1319(dataIn[1319]),
.io_parallelIn_1320(dataIn[1320]),
.io_parallelIn_1321(dataIn[1321]),
.io_parallelIn_1322(dataIn[1322]),
.io_parallelIn_1323(dataIn[1323]),
.io_parallelIn_1324(dataIn[1324]),
.io_parallelIn_1325(dataIn[1325]),
.io_parallelIn_1326(dataIn[1326]),
.io_parallelIn_1327(dataIn[1327]),
.io_parallelIn_1328(dataIn[1328]),
.io_parallelIn_1329(dataIn[1329]),
.io_parallelIn_1330(dataIn[1330]),
.io_parallelIn_1331(dataIn[1331]),
.io_parallelIn_1332(dataIn[1332]),
.io_parallelIn_1333(dataIn[1333]),
.io_parallelIn_1334(dataIn[1334]),
.io_parallelIn_1335(dataIn[1335]),
.io_parallelIn_1336(dataIn[1336]),
.io_parallelIn_1337(dataIn[1337]),
.io_parallelIn_1338(dataIn[1338]),
.io_parallelIn_1339(dataIn[1339]),
.io_parallelIn_1340(dataIn[1340]),
.io_parallelIn_1341(dataIn[1341]),
.io_parallelIn_1342(dataIn[1342]),
.io_parallelIn_1343(dataIn[1343]),
.io_parallelIn_1344(dataIn[1344]),
.io_parallelIn_1345(dataIn[1345]),
.io_parallelIn_1346(dataIn[1346]),
.io_parallelIn_1347(dataIn[1347]),
.io_parallelIn_1348(dataIn[1348]),
.io_parallelIn_1349(dataIn[1349]),
.io_parallelIn_1350(dataIn[1350]),
.io_parallelIn_1351(dataIn[1351]),
.io_parallelIn_1352(dataIn[1352]),
.io_parallelIn_1353(dataIn[1353]),
.io_parallelIn_1354(dataIn[1354]),
.io_parallelIn_1355(dataIn[1355]),
.io_parallelIn_1356(dataIn[1356]),
.io_parallelIn_1357(dataIn[1357]),
.io_parallelIn_1358(dataIn[1358]),
.io_parallelIn_1359(dataIn[1359]),
.io_parallelIn_1360(dataIn[1360]),
.io_parallelIn_1361(dataIn[1361]),
.io_parallelIn_1362(dataIn[1362]),
.io_parallelIn_1363(dataIn[1363]),
.io_parallelIn_1364(dataIn[1364]),
.io_parallelIn_1365(dataIn[1365]),
.io_parallelIn_1366(dataIn[1366]),
.io_parallelIn_1367(dataIn[1367]),
.io_parallelIn_1368(dataIn[1368]),
.io_parallelIn_1369(dataIn[1369]),
.io_parallelIn_1370(dataIn[1370]),
.io_parallelIn_1371(dataIn[1371]),
.io_parallelIn_1372(dataIn[1372]),
.io_parallelIn_1373(dataIn[1373]),
.io_parallelIn_1374(dataIn[1374]),
.io_parallelIn_1375(dataIn[1375]),
.io_parallelIn_1376(dataIn[1376]),
.io_parallelIn_1377(dataIn[1377]),
.io_parallelIn_1378(dataIn[1378]),
.io_parallelIn_1379(dataIn[1379]),
.io_parallelIn_1380(dataIn[1380]),
.io_parallelIn_1381(dataIn[1381]),
.io_parallelIn_1382(dataIn[1382]),
.io_parallelIn_1383(dataIn[1383]),
.io_parallelIn_1384(dataIn[1384]),
.io_parallelIn_1385(dataIn[1385]),
.io_parallelIn_1386(dataIn[1386]),
.io_parallelIn_1387(dataIn[1387]),
.io_parallelIn_1388(dataIn[1388]),
.io_parallelIn_1389(dataIn[1389]),
.io_parallelIn_1390(dataIn[1390]),
.io_parallelIn_1391(dataIn[1391]),
.io_parallelIn_1392(dataIn[1392]),
.io_parallelIn_1393(dataIn[1393]),
.io_parallelIn_1394(dataIn[1394]),
.io_parallelIn_1395(dataIn[1395]),
.io_parallelIn_1396(dataIn[1396]),
.io_parallelIn_1397(dataIn[1397]),
.io_parallelIn_1398(dataIn[1398]),
.io_parallelIn_1399(dataIn[1399]),
.io_parallelIn_1400(dataIn[1400]),
.io_parallelIn_1401(dataIn[1401]),
.io_parallelIn_1402(dataIn[1402]),
.io_parallelIn_1403(dataIn[1403]),
.io_parallelIn_1404(dataIn[1404]),
.io_parallelIn_1405(dataIn[1405]),
.io_parallelIn_1406(dataIn[1406]),
.io_parallelIn_1407(dataIn[1407]),
.io_parallelIn_1408(dataIn[1408]),
.io_parallelIn_1409(dataIn[1409]),
.io_parallelIn_1410(dataIn[1410]),
.io_parallelIn_1411(dataIn[1411]),
.io_parallelIn_1412(dataIn[1412]),
.io_parallelIn_1413(dataIn[1413]),
.io_parallelIn_1414(dataIn[1414]),
.io_parallelIn_1415(dataIn[1415]),
.io_parallelIn_1416(dataIn[1416]),
.io_parallelIn_1417(dataIn[1417]),
.io_parallelIn_1418(dataIn[1418]),
.io_parallelIn_1419(dataIn[1419]),
.io_parallelIn_1420(dataIn[1420]),
.io_parallelIn_1421(dataIn[1421]),
.io_parallelIn_1422(dataIn[1422]),
.io_parallelIn_1423(dataIn[1423]),
.io_parallelIn_1424(dataIn[1424]),
.io_parallelIn_1425(dataIn[1425]),
.io_parallelIn_1426(dataIn[1426]),
.io_parallelIn_1427(dataIn[1427]),
.io_parallelIn_1428(dataIn[1428]),
.io_parallelIn_1429(dataIn[1429]),
.io_parallelIn_1430(dataIn[1430]),
.io_parallelIn_1431(dataIn[1431]),
.io_parallelIn_1432(dataIn[1432]),
.io_parallelIn_1433(dataIn[1433]),
.io_parallelIn_1434(dataIn[1434]),
.io_parallelIn_1435(dataIn[1435]),
.io_parallelIn_1436(dataIn[1436]),
.io_parallelIn_1437(dataIn[1437]),
.io_parallelIn_1438(dataIn[1438]),
.io_parallelIn_1439(dataIn[1439]),
.io_parallelIn_1440(dataIn[1440]),
.io_parallelIn_1441(dataIn[1441]),
.io_parallelIn_1442(dataIn[1442]),
.io_parallelIn_1443(dataIn[1443]),
.io_parallelIn_1444(dataIn[1444]),
.io_parallelIn_1445(dataIn[1445]),
.io_parallelIn_1446(dataIn[1446]),
.io_parallelIn_1447(dataIn[1447]),
.io_parallelIn_1448(dataIn[1448]),
.io_parallelIn_1449(dataIn[1449]),
.io_parallelIn_1450(dataIn[1450]),
.io_parallelIn_1451(dataIn[1451]),
.io_parallelIn_1452(dataIn[1452]),
.io_parallelIn_1453(dataIn[1453]),
.io_parallelIn_1454(dataIn[1454]),
.io_parallelIn_1455(dataIn[1455]),
.io_parallelIn_1456(dataIn[1456]),
.io_parallelIn_1457(dataIn[1457]),
.io_parallelIn_1458(dataIn[1458]),
.io_parallelIn_1459(dataIn[1459]),
.io_parallelIn_1460(dataIn[1460]),
.io_parallelIn_1461(dataIn[1461]),
.io_parallelIn_1462(dataIn[1462]),
.io_parallelIn_1463(dataIn[1463]),
.io_parallelIn_1464(dataIn[1464]),
.io_parallelIn_1465(dataIn[1465]),
.io_parallelIn_1466(dataIn[1466]),
.io_parallelIn_1467(dataIn[1467]),
.io_parallelIn_1468(dataIn[1468]),
.io_parallelIn_1469(dataIn[1469]),
.io_parallelIn_1470(dataIn[1470]),
.io_parallelIn_1471(dataIn[1471]),
.io_parallelIn_1472(dataIn[1472]),
.io_parallelIn_1473(dataIn[1473]),
.io_parallelIn_1474(dataIn[1474]),
.io_parallelIn_1475(dataIn[1475]),
.io_parallelIn_1476(dataIn[1476]),
.io_parallelIn_1477(dataIn[1477]),
.io_parallelIn_1478(dataIn[1478]),
.io_parallelIn_1479(dataIn[1479]),
.io_parallelIn_1480(dataIn[1480]),
.io_parallelIn_1481(dataIn[1481]),
.io_parallelIn_1482(dataIn[1482]),
.io_parallelIn_1483(dataIn[1483]),
.io_parallelIn_1484(dataIn[1484]),
.io_parallelIn_1485(dataIn[1485]),
.io_parallelIn_1486(dataIn[1486]),
.io_parallelIn_1487(dataIn[1487]),
.io_parallelIn_1488(dataIn[1488]),
.io_parallelIn_1489(dataIn[1489]),
.io_parallelIn_1490(dataIn[1490]),
.io_parallelIn_1491(dataIn[1491]),
.io_parallelIn_1492(dataIn[1492]),
.io_parallelIn_1493(dataIn[1493]),
.io_parallelIn_1494(dataIn[1494]),
.io_parallelIn_1495(dataIn[1495]),
.io_parallelIn_1496(dataIn[1496]),
.io_parallelIn_1497(dataIn[1497]),
.io_parallelIn_1498(dataIn[1498]),
.io_parallelIn_1499(dataIn[1499]),
.io_parallelIn_1500(dataIn[1500]),
.io_parallelIn_1501(dataIn[1501]),
.io_parallelIn_1502(dataIn[1502]),
.io_parallelIn_1503(dataIn[1503]),
.io_parallelIn_1504(dataIn[1504]),
.io_parallelIn_1505(dataIn[1505]),
.io_parallelIn_1506(dataIn[1506]),
.io_parallelIn_1507(dataIn[1507]),
.io_parallelIn_1508(dataIn[1508]),
.io_parallelIn_1509(dataIn[1509]),
.io_parallelIn_1510(dataIn[1510]),
.io_parallelIn_1511(dataIn[1511]),
.io_parallelIn_1512(dataIn[1512]),
.io_parallelIn_1513(dataIn[1513]),
.io_parallelIn_1514(dataIn[1514]),
.io_parallelIn_1515(dataIn[1515]),
.io_parallelIn_1516(dataIn[1516]),
.io_parallelIn_1517(dataIn[1517]),
.io_parallelIn_1518(dataIn[1518]),
.io_parallelIn_1519(dataIn[1519]),
.io_parallelIn_1520(dataIn[1520]),
.io_parallelIn_1521(dataIn[1521]),
.io_parallelIn_1522(dataIn[1522]),
.io_parallelIn_1523(dataIn[1523]),
.io_parallelIn_1524(dataIn[1524]),
.io_parallelIn_1525(dataIn[1525]),
.io_parallelIn_1526(dataIn[1526]),
.io_parallelIn_1527(dataIn[1527]),
.io_parallelIn_1528(dataIn[1528]),
.io_parallelIn_1529(dataIn[1529]),
.io_parallelIn_1530(dataIn[1530]),
.io_parallelIn_1531(dataIn[1531]),
.io_parallelIn_1532(dataIn[1532]),
.io_parallelIn_1533(dataIn[1533]),
.io_parallelIn_1534(dataIn[1534]),
.io_parallelIn_1535(dataIn[1535]),
.io_parallelIn_1536(dataIn[1536]),
.io_parallelIn_1537(dataIn[1537]),
.io_parallelIn_1538(dataIn[1538]),
.io_parallelIn_1539(dataIn[1539]),
.io_parallelIn_1540(dataIn[1540]),
.io_parallelIn_1541(dataIn[1541]),
.io_parallelIn_1542(dataIn[1542]),
.io_parallelIn_1543(dataIn[1543]),
.io_parallelIn_1544(dataIn[1544]),
.io_parallelIn_1545(dataIn[1545]),
.io_parallelIn_1546(dataIn[1546]),
.io_parallelIn_1547(dataIn[1547]),
.io_parallelIn_1548(dataIn[1548]),
.io_parallelIn_1549(dataIn[1549]),
.io_parallelIn_1550(dataIn[1550]),
.io_parallelIn_1551(dataIn[1551]),
.io_parallelIn_1552(dataIn[1552]),
.io_parallelIn_1553(dataIn[1553]),
.io_parallelIn_1554(dataIn[1554]),
.io_parallelIn_1555(dataIn[1555]),
.io_parallelIn_1556(dataIn[1556]),
.io_parallelIn_1557(dataIn[1557]),
.io_parallelIn_1558(dataIn[1558]),
.io_parallelIn_1559(dataIn[1559]),
.io_parallelIn_1560(dataIn[1560]),
.io_parallelIn_1561(dataIn[1561]),
.io_parallelIn_1562(dataIn[1562]),
.io_parallelIn_1563(dataIn[1563]),
.io_parallelIn_1564(dataIn[1564]),
.io_parallelIn_1565(dataIn[1565]),
.io_parallelIn_1566(dataIn[1566]),
.io_parallelIn_1567(dataIn[1567]),
.io_parallelIn_1568(dataIn[1568]),
.io_parallelIn_1569(dataIn[1569]),
.io_parallelIn_1570(dataIn[1570]),
.io_parallelIn_1571(dataIn[1571]),
.io_parallelIn_1572(dataIn[1572]),
.io_parallelIn_1573(dataIn[1573]),
.io_parallelIn_1574(dataIn[1574]),
.io_parallelIn_1575(dataIn[1575]),
.io_parallelIn_1576(dataIn[1576]),
.io_parallelIn_1577(dataIn[1577]),
.io_parallelIn_1578(dataIn[1578]),
.io_parallelIn_1579(dataIn[1579]),
.io_parallelIn_1580(dataIn[1580]),
.io_parallelIn_1581(dataIn[1581]),
.io_parallelIn_1582(dataIn[1582]),
.io_parallelIn_1583(dataIn[1583]),
.io_parallelIn_1584(dataIn[1584]),
.io_parallelIn_1585(dataIn[1585]),
.io_parallelIn_1586(dataIn[1586]),
.io_parallelIn_1587(dataIn[1587]),
.io_parallelIn_1588(dataIn[1588]),
.io_parallelIn_1589(dataIn[1589]),
.io_parallelIn_1590(dataIn[1590]),
.io_parallelIn_1591(dataIn[1591]),
.io_parallelIn_1592(dataIn[1592]),
.io_parallelIn_1593(dataIn[1593]),
.io_parallelIn_1594(dataIn[1594]),
.io_parallelIn_1595(dataIn[1595]),
.io_parallelIn_1596(dataIn[1596]),
.io_parallelIn_1597(dataIn[1597]),
.io_parallelIn_1598(dataIn[1598]),
.io_parallelIn_1599(dataIn[1599]),
.io_parallelIn_1600(dataIn[1600]),
.io_parallelIn_1601(dataIn[1601]),
.io_parallelIn_1602(dataIn[1602]),
.io_parallelIn_1603(dataIn[1603]),
.io_parallelIn_1604(dataIn[1604]),
.io_parallelIn_1605(dataIn[1605]),
.io_parallelIn_1606(dataIn[1606]),
.io_parallelIn_1607(dataIn[1607]),
.io_parallelIn_1608(dataIn[1608]),
.io_parallelIn_1609(dataIn[1609]),
.io_parallelIn_1610(dataIn[1610]),
.io_parallelIn_1611(dataIn[1611]),
.io_parallelIn_1612(dataIn[1612]),
.io_parallelIn_1613(dataIn[1613]),
.io_parallelIn_1614(dataIn[1614]),
.io_parallelIn_1615(dataIn[1615]),
.io_parallelIn_1616(dataIn[1616]),
.io_parallelIn_1617(dataIn[1617]),
.io_parallelIn_1618(dataIn[1618]),
.io_parallelIn_1619(dataIn[1619]),
.io_parallelIn_1620(dataIn[1620]),
.io_parallelIn_1621(dataIn[1621]),
.io_parallelIn_1622(dataIn[1622]),
.io_parallelIn_1623(dataIn[1623]),
.io_parallelIn_1624(dataIn[1624]),
.io_parallelIn_1625(dataIn[1625]),
.io_parallelIn_1626(dataIn[1626]),
.io_parallelIn_1627(dataIn[1627]),
.io_parallelIn_1628(dataIn[1628]),
.io_parallelIn_1629(dataIn[1629]),
.io_parallelIn_1630(dataIn[1630]),
.io_parallelIn_1631(dataIn[1631]),
.io_parallelIn_1632(dataIn[1632]),
.io_parallelIn_1633(dataIn[1633]),
.io_parallelIn_1634(dataIn[1634]),
.io_parallelIn_1635(dataIn[1635]),
.io_parallelIn_1636(dataIn[1636]),
.io_parallelIn_1637(dataIn[1637]),
.io_parallelIn_1638(dataIn[1638]),
.io_parallelIn_1639(dataIn[1639]),
.io_parallelIn_1640(dataIn[1640]),
.io_parallelIn_1641(dataIn[1641]),
.io_parallelIn_1642(dataIn[1642]),
.io_parallelIn_1643(dataIn[1643]),
.io_parallelIn_1644(dataIn[1644]),
.io_parallelIn_1645(dataIn[1645]),
.io_parallelIn_1646(dataIn[1646]),
.io_parallelIn_1647(dataIn[1647]),
.io_parallelIn_1648(dataIn[1648]),
.io_parallelIn_1649(dataIn[1649]),
.io_parallelIn_1650(dataIn[1650]),
.io_parallelIn_1651(dataIn[1651]),
.io_parallelIn_1652(dataIn[1652]),
.io_parallelIn_1653(dataIn[1653]),
.io_parallelIn_1654(dataIn[1654]),
.io_parallelIn_1655(dataIn[1655]),
.io_parallelIn_1656(dataIn[1656]),
.io_parallelIn_1657(dataIn[1657]),
.io_parallelIn_1658(dataIn[1658]),
.io_parallelIn_1659(dataIn[1659]),
.io_parallelIn_1660(dataIn[1660]),
.io_parallelIn_1661(dataIn[1661]),
.io_parallelIn_1662(dataIn[1662]),
.io_parallelIn_1663(dataIn[1663]),
.io_parallelIn_1664(dataIn[1664]),
.io_parallelIn_1665(dataIn[1665]),
.io_parallelIn_1666(dataIn[1666]),
.io_parallelIn_1667(dataIn[1667]),
.io_parallelIn_1668(dataIn[1668]),
.io_parallelIn_1669(dataIn[1669]),
.io_parallelIn_1670(dataIn[1670]),
.io_parallelIn_1671(dataIn[1671]),
.io_parallelIn_1672(dataIn[1672]),
.io_parallelIn_1673(dataIn[1673]),
.io_parallelIn_1674(dataIn[1674]),
.io_parallelIn_1675(dataIn[1675]),
.io_parallelIn_1676(dataIn[1676]),
.io_parallelIn_1677(dataIn[1677]),
.io_parallelIn_1678(dataIn[1678]),
.io_parallelIn_1679(dataIn[1679]),
.io_parallelIn_1680(dataIn[1680]),
.io_parallelIn_1681(dataIn[1681]),
.io_parallelIn_1682(dataIn[1682]),
.io_parallelIn_1683(dataIn[1683]),
.io_parallelIn_1684(dataIn[1684]),
.io_parallelIn_1685(dataIn[1685]),
.io_parallelIn_1686(dataIn[1686]),
.io_parallelIn_1687(dataIn[1687]),
.io_parallelIn_1688(dataIn[1688]),
.io_parallelIn_1689(dataIn[1689]),
.io_parallelIn_1690(dataIn[1690]),
.io_parallelIn_1691(dataIn[1691]),
.io_parallelIn_1692(dataIn[1692]),
.io_parallelIn_1693(dataIn[1693]),
.io_parallelIn_1694(dataIn[1694]),
.io_parallelIn_1695(dataIn[1695]),
.io_parallelIn_1696(dataIn[1696]),
.io_parallelIn_1697(dataIn[1697]),
.io_parallelIn_1698(dataIn[1698]),
.io_parallelIn_1699(dataIn[1699]),
.io_parallelIn_1700(dataIn[1700]),
.io_parallelIn_1701(dataIn[1701]),
.io_parallelIn_1702(dataIn[1702]),
.io_parallelIn_1703(dataIn[1703]),
.io_parallelIn_1704(dataIn[1704]),
.io_parallelIn_1705(dataIn[1705]),
.io_parallelIn_1706(dataIn[1706]),
.io_parallelIn_1707(dataIn[1707]),
.io_parallelIn_1708(dataIn[1708]),
.io_parallelIn_1709(dataIn[1709]),
.io_parallelIn_1710(dataIn[1710]),
.io_parallelIn_1711(dataIn[1711]),
.io_parallelIn_1712(dataIn[1712]),
.io_parallelIn_1713(dataIn[1713]),
.io_parallelIn_1714(dataIn[1714]),
.io_parallelIn_1715(dataIn[1715]),
.io_parallelIn_1716(dataIn[1716]),
.io_parallelIn_1717(dataIn[1717]),
.io_parallelIn_1718(dataIn[1718]),
.io_parallelIn_1719(dataIn[1719]),
.io_parallelIn_1720(dataIn[1720]),
.io_parallelIn_1721(dataIn[1721]),
.io_parallelIn_1722(dataIn[1722]),
.io_parallelIn_1723(dataIn[1723]),
.io_parallelIn_1724(dataIn[1724]),
.io_parallelIn_1725(dataIn[1725]),
.io_parallelIn_1726(dataIn[1726]),
.io_parallelIn_1727(dataIn[1727]),
.io_parallelIn_1728(dataIn[1728]),
.io_parallelIn_1729(dataIn[1729]),
.io_parallelIn_1730(dataIn[1730]),
.io_parallelIn_1731(dataIn[1731]),
.io_parallelIn_1732(dataIn[1732]),
.io_parallelIn_1733(dataIn[1733]),
.io_parallelIn_1734(dataIn[1734]),
.io_parallelIn_1735(dataIn[1735]),
.io_parallelIn_1736(dataIn[1736]),
.io_parallelIn_1737(dataIn[1737]),
.io_parallelIn_1738(dataIn[1738]),
.io_parallelIn_1739(dataIn[1739]),
.io_parallelIn_1740(dataIn[1740]),
.io_parallelIn_1741(dataIn[1741]),
.io_parallelIn_1742(dataIn[1742]),
.io_parallelIn_1743(dataIn[1743]),
.io_parallelIn_1744(dataIn[1744]),
.io_parallelIn_1745(dataIn[1745]),
.io_parallelIn_1746(dataIn[1746]),
.io_parallelIn_1747(dataIn[1747]),
.io_parallelIn_1748(dataIn[1748]),
.io_parallelIn_1749(dataIn[1749]),
.io_parallelIn_1750(dataIn[1750]),
.io_parallelIn_1751(dataIn[1751]),
.io_parallelIn_1752(dataIn[1752]),
.io_parallelIn_1753(dataIn[1753]),
.io_parallelIn_1754(dataIn[1754]),
.io_parallelIn_1755(dataIn[1755]),
.io_parallelIn_1756(dataIn[1756]),
.io_parallelIn_1757(dataIn[1757]),
.io_parallelIn_1758(dataIn[1758]),
.io_parallelIn_1759(dataIn[1759]),
.io_parallelIn_1760(dataIn[1760]),
.io_parallelIn_1761(dataIn[1761]),
.io_parallelIn_1762(dataIn[1762]),
.io_parallelIn_1763(dataIn[1763]),
.io_parallelIn_1764(dataIn[1764]),
.io_parallelIn_1765(dataIn[1765]),
.io_parallelIn_1766(dataIn[1766]),
.io_parallelIn_1767(dataIn[1767]),
.io_parallelIn_1768(dataIn[1768]),
.io_parallelIn_1769(dataIn[1769]),
.io_parallelIn_1770(dataIn[1770]),
.io_parallelIn_1771(dataIn[1771]),
.io_parallelIn_1772(dataIn[1772]),
.io_parallelIn_1773(dataIn[1773]),
.io_parallelIn_1774(dataIn[1774]),
.io_parallelIn_1775(dataIn[1775]),
.io_parallelIn_1776(dataIn[1776]),
.io_parallelIn_1777(dataIn[1777]),
.io_parallelIn_1778(dataIn[1778]),
.io_parallelIn_1779(dataIn[1779]),
.io_parallelIn_1780(dataIn[1780]),
.io_parallelIn_1781(dataIn[1781]),
.io_parallelIn_1782(dataIn[1782]),
.io_parallelIn_1783(dataIn[1783]),
.io_parallelIn_1784(dataIn[1784]),
.io_parallelIn_1785(dataIn[1785]),
.io_parallelIn_1786(dataIn[1786]),
.io_parallelIn_1787(dataIn[1787]),
.io_parallelIn_1788(dataIn[1788]),
.io_parallelIn_1789(dataIn[1789]),
.io_parallelIn_1790(dataIn[1790]),
.io_parallelIn_1791(dataIn[1791]),
.io_parallelIn_1792(dataIn[1792]),
.io_parallelIn_1793(dataIn[1793]),
.io_parallelIn_1794(dataIn[1794]),
.io_parallelIn_1795(dataIn[1795]),
.io_parallelIn_1796(dataIn[1796]),
.io_parallelIn_1797(dataIn[1797]),
.io_parallelIn_1798(dataIn[1798]),
.io_parallelIn_1799(dataIn[1799]),
.io_parallelIn_1800(dataIn[1800]),
.io_parallelIn_1801(dataIn[1801]),
.io_parallelIn_1802(dataIn[1802]),
.io_parallelIn_1803(dataIn[1803]),
.io_parallelIn_1804(dataIn[1804]),
.io_parallelIn_1805(dataIn[1805]),
.io_parallelIn_1806(dataIn[1806]),
.io_parallelIn_1807(dataIn[1807]),
.io_parallelIn_1808(dataIn[1808]),
.io_parallelIn_1809(dataIn[1809]),
.io_parallelIn_1810(dataIn[1810]),
.io_parallelIn_1811(dataIn[1811]),
.io_parallelIn_1812(dataIn[1812]),
.io_parallelIn_1813(dataIn[1813]),
.io_parallelIn_1814(dataIn[1814]),
.io_parallelIn_1815(dataIn[1815]),
.io_parallelIn_1816(dataIn[1816]),
.io_parallelIn_1817(dataIn[1817]),
.io_parallelIn_1818(dataIn[1818]),
.io_parallelIn_1819(dataIn[1819]),
.io_parallelIn_1820(dataIn[1820]),
.io_parallelIn_1821(dataIn[1821]),
.io_parallelIn_1822(dataIn[1822]),
.io_parallelIn_1823(dataIn[1823]),
.io_parallelIn_1824(dataIn[1824]),
.io_parallelIn_1825(dataIn[1825]),
.io_parallelIn_1826(dataIn[1826]),
.io_parallelIn_1827(dataIn[1827]),
.io_parallelIn_1828(dataIn[1828]),
.io_parallelIn_1829(dataIn[1829]),
.io_parallelIn_1830(dataIn[1830]),
.io_parallelIn_1831(dataIn[1831]),
.io_parallelIn_1832(dataIn[1832]),
.io_parallelIn_1833(dataIn[1833]),
.io_parallelIn_1834(dataIn[1834]),
.io_parallelIn_1835(dataIn[1835]),
.io_parallelIn_1836(dataIn[1836]),
.io_parallelIn_1837(dataIn[1837]),
.io_parallelIn_1838(dataIn[1838]),
.io_parallelIn_1839(dataIn[1839]),
.io_parallelIn_1840(dataIn[1840]),
.io_parallelIn_1841(dataIn[1841]),
.io_parallelIn_1842(dataIn[1842]),
.io_parallelIn_1843(dataIn[1843]),
.io_parallelIn_1844(dataIn[1844]),
.io_parallelIn_1845(dataIn[1845]),
.io_parallelIn_1846(dataIn[1846]),
.io_parallelIn_1847(dataIn[1847]),
.io_parallelIn_1848(dataIn[1848]),
.io_parallelIn_1849(dataIn[1849]),
.io_parallelIn_1850(dataIn[1850]),
.io_parallelIn_1851(dataIn[1851]),
.io_parallelIn_1852(dataIn[1852]),
.io_parallelIn_1853(dataIn[1853]),
.io_parallelIn_1854(dataIn[1854]),
.io_parallelIn_1855(dataIn[1855]),
.io_parallelIn_1856(dataIn[1856]),
.io_parallelIn_1857(dataIn[1857]),
.io_parallelIn_1858(dataIn[1858]),
.io_parallelIn_1859(dataIn[1859]),
.io_parallelIn_1860(dataIn[1860]),
.io_parallelIn_1861(dataIn[1861]),
.io_parallelIn_1862(dataIn[1862]),
.io_parallelIn_1863(dataIn[1863]),
.io_parallelIn_1864(dataIn[1864]),
.io_parallelIn_1865(dataIn[1865]),
.io_parallelIn_1866(dataIn[1866]),
.io_parallelIn_1867(dataIn[1867]),
.io_parallelIn_1868(dataIn[1868]),
.io_parallelIn_1869(dataIn[1869]),
.io_parallelIn_1870(dataIn[1870]),
.io_parallelIn_1871(dataIn[1871]),
.io_parallelIn_1872(dataIn[1872]),
.io_parallelIn_1873(dataIn[1873]),
.io_parallelIn_1874(dataIn[1874]),
.io_parallelIn_1875(dataIn[1875]),
.io_parallelIn_1876(dataIn[1876]),
.io_parallelIn_1877(dataIn[1877]),
.io_parallelIn_1878(dataIn[1878]),
.io_parallelIn_1879(dataIn[1879]),
.io_parallelIn_1880(dataIn[1880]),
.io_parallelIn_1881(dataIn[1881]),
.io_parallelIn_1882(dataIn[1882]),
.io_parallelIn_1883(dataIn[1883]),
.io_parallelIn_1884(dataIn[1884]),
.io_parallelIn_1885(dataIn[1885]),
.io_parallelIn_1886(dataIn[1886]),
.io_parallelIn_1887(dataIn[1887]),
.io_parallelIn_1888(dataIn[1888]),
.io_parallelIn_1889(dataIn[1889]),
.io_parallelIn_1890(dataIn[1890]),
.io_parallelIn_1891(dataIn[1891]),
.io_parallelIn_1892(dataIn[1892]),
.io_parallelIn_1893(dataIn[1893]),
.io_parallelIn_1894(dataIn[1894]),
.io_parallelIn_1895(dataIn[1895]),
.io_parallelIn_1896(dataIn[1896]),
.io_parallelIn_1897(dataIn[1897]),
.io_parallelIn_1898(dataIn[1898]),
.io_parallelIn_1899(dataIn[1899]),
.io_parallelIn_1900(dataIn[1900]),
.io_parallelIn_1901(dataIn[1901]),
.io_parallelIn_1902(dataIn[1902]),
.io_parallelIn_1903(dataIn[1903]),
.io_parallelIn_1904(dataIn[1904]),
.io_parallelIn_1905(dataIn[1905]),
.io_parallelIn_1906(dataIn[1906]),
.io_parallelIn_1907(dataIn[1907]),
.io_parallelIn_1908(dataIn[1908]),
.io_parallelIn_1909(dataIn[1909]),
.io_parallelIn_1910(dataIn[1910]),
.io_parallelIn_1911(dataIn[1911]),
.io_parallelIn_1912(dataIn[1912]),
.io_parallelIn_1913(dataIn[1913]),
.io_parallelIn_1914(dataIn[1914]),
.io_parallelIn_1915(dataIn[1915]),
.io_parallelIn_1916(dataIn[1916]),
.io_parallelIn_1917(dataIn[1917]),
.io_parallelIn_1918(dataIn[1918]),
.io_parallelIn_1919(dataIn[1919]),
.io_parallelIn_1920(dataIn[1920]),
.io_parallelIn_1921(dataIn[1921]),
.io_parallelIn_1922(dataIn[1922]),
.io_parallelIn_1923(dataIn[1923]),
.io_parallelIn_1924(dataIn[1924]),
.io_parallelIn_1925(dataIn[1925]),
.io_parallelIn_1926(dataIn[1926]),
.io_parallelIn_1927(dataIn[1927]),
.io_parallelIn_1928(dataIn[1928]),
.io_parallelIn_1929(dataIn[1929]),
.io_parallelIn_1930(dataIn[1930]),
.io_parallelIn_1931(dataIn[1931]),
.io_parallelIn_1932(dataIn[1932]),
.io_parallelIn_1933(dataIn[1933]),
.io_parallelIn_1934(dataIn[1934]),
.io_parallelIn_1935(dataIn[1935]),
.io_parallelIn_1936(dataIn[1936]),
.io_parallelIn_1937(dataIn[1937]),
.io_parallelIn_1938(dataIn[1938]),
.io_parallelIn_1939(dataIn[1939]),
.io_parallelIn_1940(dataIn[1940]),
.io_parallelIn_1941(dataIn[1941]),
.io_parallelIn_1942(dataIn[1942]),
.io_parallelIn_1943(dataIn[1943]),
.io_parallelIn_1944(dataIn[1944]),
.io_parallelIn_1945(dataIn[1945]),
.io_parallelIn_1946(dataIn[1946]),
.io_parallelIn_1947(dataIn[1947]),
.io_parallelIn_1948(dataIn[1948]),
.io_parallelIn_1949(dataIn[1949]),
.io_parallelIn_1950(dataIn[1950]),
.io_parallelIn_1951(dataIn[1951]),
.io_parallelIn_1952(dataIn[1952]),
.io_parallelIn_1953(dataIn[1953]),
.io_parallelIn_1954(dataIn[1954]),
.io_parallelIn_1955(dataIn[1955]),
.io_parallelIn_1956(dataIn[1956]),
.io_parallelIn_1957(dataIn[1957]),
.io_parallelIn_1958(dataIn[1958]),
.io_parallelIn_1959(dataIn[1959]),
.io_parallelIn_1960(dataIn[1960]),
.io_parallelIn_1961(dataIn[1961]),
.io_parallelIn_1962(dataIn[1962]),
.io_parallelIn_1963(dataIn[1963]),
.io_parallelIn_1964(dataIn[1964]),
.io_parallelIn_1965(dataIn[1965]),
.io_parallelIn_1966(dataIn[1966]),
.io_parallelIn_1967(dataIn[1967]),
.io_parallelIn_1968(dataIn[1968]),
.io_parallelIn_1969(dataIn[1969]),
.io_parallelIn_1970(dataIn[1970]),
.io_parallelIn_1971(dataIn[1971]),
.io_parallelIn_1972(dataIn[1972]),
.io_parallelIn_1973(dataIn[1973]),
.io_parallelIn_1974(dataIn[1974]),
.io_parallelIn_1975(dataIn[1975]),
.io_parallelIn_1976(dataIn[1976]),
.io_parallelIn_1977(dataIn[1977]),
.io_parallelIn_1978(dataIn[1978]),
.io_parallelIn_1979(dataIn[1979]),
.io_parallelIn_1980(dataIn[1980]),
.io_parallelIn_1981(dataIn[1981]),
.io_parallelIn_1982(dataIn[1982]),
.io_parallelIn_1983(dataIn[1983]),
.io_parallelIn_1984(dataIn[1984]),
.io_parallelIn_1985(dataIn[1985]),
.io_parallelIn_1986(dataIn[1986]),
.io_parallelIn_1987(dataIn[1987]),
.io_parallelIn_1988(dataIn[1988]),
.io_parallelIn_1989(dataIn[1989]),
.io_parallelIn_1990(dataIn[1990]),
.io_parallelIn_1991(dataIn[1991]),
.io_parallelIn_1992(dataIn[1992]),
.io_parallelIn_1993(dataIn[1993]),
.io_parallelIn_1994(dataIn[1994]),
.io_parallelIn_1995(dataIn[1995]),
.io_parallelIn_1996(dataIn[1996]),
.io_parallelIn_1997(dataIn[1997]),
.io_parallelIn_1998(dataIn[1998]),
.io_parallelIn_1999(dataIn[1999]),
.io_parallelIn_2000(dataIn[2000]),
.io_parallelIn_2001(dataIn[2001]),
.io_parallelIn_2002(dataIn[2002]),
.io_parallelIn_2003(dataIn[2003]),
.io_parallelIn_2004(dataIn[2004]),
.io_parallelIn_2005(dataIn[2005]),
.io_parallelIn_2006(dataIn[2006]),
.io_parallelIn_2007(dataIn[2007]),
.io_parallelIn_2008(dataIn[2008]),
.io_parallelIn_2009(dataIn[2009]),
.io_parallelIn_2010(dataIn[2010]),
.io_parallelIn_2011(dataIn[2011]),
.io_parallelIn_2012(dataIn[2012]),
.io_parallelIn_2013(dataIn[2013]),
.io_parallelIn_2014(dataIn[2014]),
.io_parallelIn_2015(dataIn[2015]),
.io_parallelIn_2016(dataIn[2016]),
.io_parallelIn_2017(dataIn[2017]),
.io_parallelIn_2018(dataIn[2018]),
.io_parallelIn_2019(dataIn[2019]),
.io_parallelIn_2020(dataIn[2020]),
.io_parallelIn_2021(dataIn[2021]),
.io_parallelIn_2022(dataIn[2022]),
.io_parallelIn_2023(dataIn[2023]),
.io_parallelIn_2024(dataIn[2024]),
.io_parallelIn_2025(dataIn[2025]),
.io_parallelIn_2026(dataIn[2026]),
.io_parallelIn_2027(dataIn[2027]),
.io_parallelIn_2028(dataIn[2028]),
.io_parallelIn_2029(dataIn[2029]),
.io_parallelIn_2030(dataIn[2030]),
.io_parallelIn_2031(dataIn[2031]),
.io_parallelIn_2032(dataIn[2032]),
.io_parallelIn_2033(dataIn[2033]),
.io_parallelIn_2034(dataIn[2034]),
.io_parallelIn_2035(dataIn[2035]),
.io_parallelIn_2036(dataIn[2036]),
.io_parallelIn_2037(dataIn[2037]),
.io_parallelIn_2038(dataIn[2038]),
.io_parallelIn_2039(dataIn[2039]),
.io_parallelIn_2040(dataIn[2040]),
.io_parallelIn_2041(dataIn[2041]),
.io_parallelIn_2042(dataIn[2042]),
.io_parallelIn_2043(dataIn[2043]),
.io_parallelIn_2044(dataIn[2044]),
.io_parallelIn_2045(dataIn[2045]),
.io_parallelIn_2046(dataIn[2046]),
.io_parallelIn_2047(dataIn[2047]),
.io_parallelIn_2048(dataIn[2048]),
.io_parallelIn_2049(dataIn[2049]),
.io_parallelIn_2050(dataIn[2050]),
.io_parallelIn_2051(dataIn[2051]),
.io_parallelIn_2052(dataIn[2052]),
.io_parallelIn_2053(dataIn[2053]),
.io_parallelIn_2054(dataIn[2054]),
.io_parallelIn_2055(dataIn[2055]),
.io_parallelIn_2056(dataIn[2056]),
.io_parallelIn_2057(dataIn[2057]),
.io_parallelIn_2058(dataIn[2058]),
.io_parallelIn_2059(dataIn[2059]),
.io_parallelIn_2060(dataIn[2060]),
.io_parallelIn_2061(dataIn[2061]),
.io_parallelIn_2062(dataIn[2062]),
.io_parallelIn_2063(dataIn[2063]),
.io_parallelIn_2064(dataIn[2064]),
.io_parallelIn_2065(dataIn[2065]),
.io_parallelIn_2066(dataIn[2066]),
.io_parallelIn_2067(dataIn[2067]),
.io_parallelIn_2068(dataIn[2068]),
.io_parallelIn_2069(dataIn[2069]),
.io_parallelIn_2070(dataIn[2070]),
.io_parallelIn_2071(dataIn[2071]),
.io_parallelIn_2072(dataIn[2072]),
.io_parallelIn_2073(dataIn[2073]),
.io_parallelIn_2074(dataIn[2074]),
.io_parallelIn_2075(dataIn[2075]),
.io_parallelIn_2076(dataIn[2076]),
.io_parallelIn_2077(dataIn[2077]),
.io_parallelIn_2078(dataIn[2078]),
.io_parallelIn_2079(dataIn[2079]),
.io_parallelIn_2080(dataIn[2080]),
.io_parallelIn_2081(dataIn[2081]),
.io_parallelIn_2082(dataIn[2082]),
.io_parallelIn_2083(dataIn[2083]),
.io_parallelIn_2084(dataIn[2084]),
.io_parallelIn_2085(dataIn[2085]),
.io_parallelIn_2086(dataIn[2086]),
.io_parallelIn_2087(dataIn[2087]),
.io_parallelIn_2088(dataIn[2088]),
.io_parallelIn_2089(dataIn[2089]),
.io_parallelIn_2090(dataIn[2090]),
.io_parallelIn_2091(dataIn[2091]),
.io_parallelIn_2092(dataIn[2092]),
.io_parallelIn_2093(dataIn[2093]),
.io_parallelIn_2094(dataIn[2094]),
.io_parallelIn_2095(dataIn[2095]),
.io_parallelIn_2096(dataIn[2096]),
.io_parallelIn_2097(dataIn[2097]),
.io_parallelIn_2098(dataIn[2098]),
.io_parallelIn_2099(dataIn[2099]),
.io_parallelIn_2100(dataIn[2100]),
.io_parallelIn_2101(dataIn[2101]),
.io_parallelIn_2102(dataIn[2102]),
.io_parallelIn_2103(dataIn[2103]),
.io_parallelIn_2104(dataIn[2104]),
.io_parallelIn_2105(dataIn[2105]),
.io_parallelIn_2106(dataIn[2106]),
.io_parallelIn_2107(dataIn[2107]),
.io_parallelIn_2108(dataIn[2108]),
.io_parallelIn_2109(dataIn[2109]),
.io_parallelIn_2110(dataIn[2110]),
.io_parallelIn_2111(dataIn[2111]),
.io_parallelIn_2112(dataIn[2112]),
.io_parallelIn_2113(dataIn[2113]),
.io_parallelIn_2114(dataIn[2114]),
.io_parallelIn_2115(dataIn[2115]),
.io_parallelIn_2116(dataIn[2116]),
.io_parallelIn_2117(dataIn[2117]),
.io_parallelIn_2118(dataIn[2118]),
.io_parallelIn_2119(dataIn[2119]),
.io_parallelIn_2120(dataIn[2120]),
.io_parallelIn_2121(dataIn[2121]),
.io_parallelIn_2122(dataIn[2122]),
.io_parallelIn_2123(dataIn[2123]),
.io_parallelIn_2124(dataIn[2124]),
.io_parallelIn_2125(dataIn[2125]),
.io_parallelIn_2126(dataIn[2126]),
.io_parallelIn_2127(dataIn[2127]),
.io_parallelIn_2128(dataIn[2128]),
.io_parallelIn_2129(dataIn[2129]),
.io_parallelIn_2130(dataIn[2130]),
.io_parallelIn_2131(dataIn[2131]),
.io_parallelIn_2132(dataIn[2132]),
.io_parallelIn_2133(dataIn[2133]),
.io_parallelIn_2134(dataIn[2134]),
.io_parallelIn_2135(dataIn[2135]),
.io_parallelIn_2136(dataIn[2136]),
.io_parallelIn_2137(dataIn[2137]),
.io_parallelIn_2138(dataIn[2138]),
.io_parallelIn_2139(dataIn[2139]),
.io_parallelIn_2140(dataIn[2140]),
.io_parallelIn_2141(dataIn[2141]),
.io_parallelIn_2142(dataIn[2142]),
.io_parallelIn_2143(dataIn[2143]),
.io_parallelIn_2144(dataIn[2144]),
.io_parallelIn_2145(dataIn[2145]),
.io_parallelIn_2146(dataIn[2146]),
.io_parallelIn_2147(dataIn[2147]),
.io_parallelIn_2148(dataIn[2148]),
.io_parallelIn_2149(dataIn[2149]),
.io_parallelIn_2150(dataIn[2150]),
.io_parallelIn_2151(dataIn[2151]),
.io_parallelIn_2152(dataIn[2152]),
.io_parallelIn_2153(dataIn[2153]),
.io_parallelIn_2154(dataIn[2154]),
.io_parallelIn_2155(dataIn[2155]),
.io_parallelIn_2156(dataIn[2156]),
.io_parallelIn_2157(dataIn[2157]),
.io_parallelIn_2158(dataIn[2158]),
.io_parallelIn_2159(dataIn[2159]),
.io_parallelIn_2160(dataIn[2160]),
.io_parallelIn_2161(dataIn[2161]),
.io_parallelIn_2162(dataIn[2162]),
.io_parallelIn_2163(dataIn[2163]),
.io_parallelIn_2164(dataIn[2164]),
.io_parallelIn_2165(dataIn[2165]),
.io_parallelIn_2166(dataIn[2166]),
.io_parallelIn_2167(dataIn[2167]),
.io_parallelIn_2168(dataIn[2168]),
.io_parallelIn_2169(dataIn[2169]),
.io_parallelIn_2170(dataIn[2170]),
.io_parallelIn_2171(dataIn[2171]),
.io_parallelIn_2172(dataIn[2172]),
.io_parallelIn_2173(dataIn[2173]),
.io_parallelIn_2174(dataIn[2174]),
.io_parallelIn_2175(dataIn[2175]),
.io_parallelIn_2176(dataIn[2176]),
.io_parallelIn_2177(dataIn[2177]),
.io_parallelIn_2178(dataIn[2178]),
.io_parallelIn_2179(dataIn[2179]),
.io_parallelIn_2180(dataIn[2180]),
.io_parallelIn_2181(dataIn[2181]),
.io_parallelIn_2182(dataIn[2182]),
.io_parallelIn_2183(dataIn[2183]),
.io_parallelIn_2184(dataIn[2184]),
.io_parallelIn_2185(dataIn[2185]),
.io_parallelIn_2186(dataIn[2186]),
.io_parallelIn_2187(dataIn[2187]),
.io_parallelIn_2188(dataIn[2188]),
.io_parallelIn_2189(dataIn[2189]),
.io_parallelIn_2190(dataIn[2190]),
.io_parallelIn_2191(dataIn[2191]),
.io_parallelIn_2192(dataIn[2192]),
.io_parallelIn_2193(dataIn[2193]),
.io_parallelIn_2194(dataIn[2194]),
.io_parallelIn_2195(dataIn[2195]),
.io_parallelIn_2196(dataIn[2196]),
.io_parallelIn_2197(dataIn[2197]),
.io_parallelIn_2198(dataIn[2198]),
.io_parallelIn_2199(dataIn[2199]),
.io_parallelIn_2200(dataIn[2200]),
.io_parallelIn_2201(dataIn[2201]),
.io_parallelIn_2202(dataIn[2202]),
.io_parallelIn_2203(dataIn[2203]),
.io_parallelIn_2204(dataIn[2204]),
.io_parallelIn_2205(dataIn[2205]),
.io_parallelIn_2206(dataIn[2206]),
.io_parallelIn_2207(dataIn[2207]),
.io_parallelIn_2208(dataIn[2208]),
.io_parallelIn_2209(dataIn[2209]),
.io_parallelIn_2210(dataIn[2210]),
.io_parallelIn_2211(dataIn[2211]),
.io_parallelIn_2212(dataIn[2212]),
.io_parallelIn_2213(dataIn[2213]),
.io_parallelIn_2214(dataIn[2214]),
.io_parallelIn_2215(dataIn[2215]),
.io_parallelIn_2216(dataIn[2216]),
.io_parallelIn_2217(dataIn[2217]),
.io_parallelIn_2218(dataIn[2218]),
.io_parallelIn_2219(dataIn[2219]),
.io_parallelIn_2220(dataIn[2220]),
.io_parallelIn_2221(dataIn[2221]),
.io_parallelIn_2222(dataIn[2222]),
.io_parallelIn_2223(dataIn[2223]),
.io_parallelIn_2224(dataIn[2224]),
.io_parallelIn_2225(dataIn[2225]),
.io_parallelIn_2226(dataIn[2226]),
.io_parallelIn_2227(dataIn[2227]),
.io_parallelIn_2228(dataIn[2228]),
.io_parallelIn_2229(dataIn[2229]),
.io_parallelIn_2230(dataIn[2230]),
.io_parallelIn_2231(dataIn[2231]),
.io_parallelIn_2232(dataIn[2232]),
.io_parallelIn_2233(dataIn[2233]),
.io_parallelIn_2234(dataIn[2234]),
.io_parallelIn_2235(dataIn[2235]),
.io_parallelIn_2236(dataIn[2236]),
.io_parallelIn_2237(dataIn[2237]),
.io_parallelIn_2238(dataIn[2238]),
.io_parallelIn_2239(dataIn[2239]),
.io_parallelIn_2240(dataIn[2240]),
.io_parallelIn_2241(dataIn[2241]),
.io_parallelIn_2242(dataIn[2242]),
.io_parallelIn_2243(dataIn[2243]),
.io_parallelIn_2244(dataIn[2244]),
.io_parallelIn_2245(dataIn[2245]),
.io_parallelIn_2246(dataIn[2246]),
.io_parallelIn_2247(dataIn[2247]),
.io_parallelIn_2248(dataIn[2248]),
.io_parallelIn_2249(dataIn[2249]),
.io_parallelIn_2250(dataIn[2250]),
.io_parallelIn_2251(dataIn[2251]),
.io_parallelIn_2252(dataIn[2252]),
.io_parallelIn_2253(dataIn[2253]),
.io_parallelIn_2254(dataIn[2254]),
.io_parallelIn_2255(dataIn[2255]),
.io_parallelIn_2256(dataIn[2256]),
.io_parallelIn_2257(dataIn[2257]),
.io_parallelIn_2258(dataIn[2258]),
.io_parallelIn_2259(dataIn[2259]),
.io_parallelIn_2260(dataIn[2260]),
.io_parallelIn_2261(dataIn[2261]),
.io_parallelIn_2262(dataIn[2262]),
.io_parallelIn_2263(dataIn[2263]),
.io_parallelIn_2264(dataIn[2264]),
.io_parallelIn_2265(dataIn[2265]),
.io_parallelIn_2266(dataIn[2266]),
.io_parallelIn_2267(dataIn[2267]),
.io_parallelIn_2268(dataIn[2268]),
.io_parallelIn_2269(dataIn[2269]),
.io_parallelIn_2270(dataIn[2270]),
.io_parallelIn_2271(dataIn[2271]),
.io_parallelIn_2272(dataIn[2272]),
.io_parallelIn_2273(dataIn[2273]),
.io_parallelIn_2274(dataIn[2274]),
.io_parallelIn_2275(dataIn[2275]),
.io_parallelIn_2276(dataIn[2276]),
.io_parallelIn_2277(dataIn[2277]),
.io_parallelIn_2278(dataIn[2278]),
.io_parallelIn_2279(dataIn[2279]),
.io_parallelIn_2280(dataIn[2280]),
.io_parallelIn_2281(dataIn[2281]),
.io_parallelIn_2282(dataIn[2282]),
.io_parallelIn_2283(dataIn[2283]),
.io_parallelIn_2284(dataIn[2284]),
.io_parallelIn_2285(dataIn[2285]),
.io_parallelIn_2286(dataIn[2286]),
.io_parallelIn_2287(dataIn[2287]),
.io_parallelIn_2288(dataIn[2288]),
.io_parallelIn_2289(dataIn[2289]),
.io_parallelIn_2290(dataIn[2290]),
.io_parallelIn_2291(dataIn[2291]),
.io_parallelIn_2292(dataIn[2292]),
.io_parallelIn_2293(dataIn[2293]),
.io_parallelIn_2294(dataIn[2294]),
.io_parallelIn_2295(dataIn[2295]),
.io_parallelIn_2296(dataIn[2296]),
.io_parallelIn_2297(dataIn[2297]),
.io_parallelIn_2298(dataIn[2298]),
.io_parallelIn_2299(dataIn[2299]),
.io_parallelIn_2300(dataIn[2300]),
.io_parallelIn_2301(dataIn[2301]),
.io_parallelIn_2302(dataIn[2302]),
.io_parallelIn_2303(dataIn[2303]),
.io_parallelIn_2304(dataIn[2304]),
.io_parallelIn_2305(dataIn[2305]),
.io_parallelIn_2306(dataIn[2306]),
.io_parallelIn_2307(dataIn[2307]),
.io_parallelIn_2308(dataIn[2308]),
.io_parallelIn_2309(dataIn[2309]),
.io_parallelIn_2310(dataIn[2310]),
.io_parallelIn_2311(dataIn[2311]),
.io_parallelIn_2312(dataIn[2312]),
.io_parallelIn_2313(dataIn[2313]),
.io_parallelIn_2314(dataIn[2314]),
.io_parallelIn_2315(dataIn[2315]),
.io_parallelIn_2316(dataIn[2316]),
.io_parallelIn_2317(dataIn[2317]),
.io_parallelIn_2318(dataIn[2318]),
.io_parallelIn_2319(dataIn[2319]),
.io_parallelIn_2320(dataIn[2320]),
.io_parallelIn_2321(dataIn[2321]),
.io_parallelIn_2322(dataIn[2322]),
.io_parallelIn_2323(dataIn[2323]),
.io_parallelIn_2324(dataIn[2324]),
.io_parallelIn_2325(dataIn[2325]),
.io_parallelIn_2326(dataIn[2326]),
.io_parallelIn_2327(dataIn[2327]),
.io_parallelIn_2328(dataIn[2328]),
.io_parallelIn_2329(dataIn[2329]),
.io_parallelIn_2330(dataIn[2330]),
.io_parallelIn_2331(dataIn[2331]),
.io_parallelIn_2332(dataIn[2332]),
.io_parallelIn_2333(dataIn[2333]),
.io_parallelIn_2334(dataIn[2334]),
.io_parallelIn_2335(dataIn[2335]),
.io_parallelIn_2336(dataIn[2336]),
.io_parallelIn_2337(dataIn[2337]),
.io_parallelIn_2338(dataIn[2338]),
.io_parallelIn_2339(dataIn[2339]),
.io_parallelIn_2340(dataIn[2340]),
.io_parallelIn_2341(dataIn[2341]),
.io_parallelIn_2342(dataIn[2342]),
.io_parallelIn_2343(dataIn[2343]),
.io_parallelIn_2344(dataIn[2344]),
.io_parallelIn_2345(dataIn[2345]),
.io_parallelIn_2346(dataIn[2346]),
.io_parallelIn_2347(dataIn[2347]),
.io_parallelIn_2348(dataIn[2348]),
.io_parallelIn_2349(dataIn[2349]),
.io_parallelIn_2350(dataIn[2350]),
.io_parallelIn_2351(dataIn[2351]),
.io_parallelIn_2352(dataIn[2352]),
.io_parallelIn_2353(dataIn[2353]),
.io_parallelIn_2354(dataIn[2354]),
.io_parallelIn_2355(dataIn[2355]),
.io_parallelIn_2356(dataIn[2356]),
.io_parallelIn_2357(dataIn[2357]),
.io_parallelIn_2358(dataIn[2358]),
.io_parallelIn_2359(dataIn[2359]),
.io_parallelIn_2360(dataIn[2360]),
.io_parallelIn_2361(dataIn[2361]),
.io_parallelIn_2362(dataIn[2362]),
.io_parallelIn_2363(dataIn[2363]),
.io_parallelIn_2364(dataIn[2364]),
.io_parallelIn_2365(dataIn[2365]),
.io_parallelIn_2366(dataIn[2366]),
.io_parallelIn_2367(dataIn[2367]),
.io_parallelIn_2368(dataIn[2368]),
.io_parallelIn_2369(dataIn[2369]),
.io_parallelIn_2370(dataIn[2370]),
.io_parallelIn_2371(dataIn[2371]),
.io_parallelIn_2372(dataIn[2372]),
.io_parallelIn_2373(dataIn[2373]),
.io_parallelIn_2374(dataIn[2374]),
.io_parallelIn_2375(dataIn[2375]),
.io_parallelIn_2376(dataIn[2376]),
.io_parallelIn_2377(dataIn[2377]),
.io_parallelIn_2378(dataIn[2378]),
.io_parallelIn_2379(dataIn[2379]),
.io_parallelIn_2380(dataIn[2380]),
.io_parallelIn_2381(dataIn[2381]),
.io_parallelIn_2382(dataIn[2382]),
.io_parallelIn_2383(dataIn[2383]),
.io_parallelIn_2384(dataIn[2384]),
.io_parallelIn_2385(dataIn[2385]),
.io_parallelIn_2386(dataIn[2386]),
.io_parallelIn_2387(dataIn[2387]),
.io_parallelIn_2388(dataIn[2388]),
.io_parallelIn_2389(dataIn[2389]),
.io_parallelIn_2390(dataIn[2390]),
.io_parallelIn_2391(dataIn[2391]),
.io_parallelIn_2392(dataIn[2392]),
.io_parallelIn_2393(dataIn[2393]),
.io_parallelIn_2394(dataIn[2394]),
.io_parallelIn_2395(dataIn[2395]),
.io_parallelIn_2396(dataIn[2396]),
.io_parallelIn_2397(dataIn[2397]),
.io_parallelIn_2398(dataIn[2398]),
.io_parallelIn_2399(dataIn[2399]),
.io_parallelIn_2400(dataIn[2400]),
.io_parallelIn_2401(dataIn[2401]),
.io_parallelIn_2402(dataIn[2402]),
.io_parallelIn_2403(dataIn[2403]),
.io_parallelIn_2404(dataIn[2404]),
.io_parallelIn_2405(dataIn[2405]),
.io_parallelIn_2406(dataIn[2406]),
.io_parallelIn_2407(dataIn[2407]),
.io_parallelIn_2408(dataIn[2408]),
.io_parallelIn_2409(dataIn[2409]),
.io_parallelIn_2410(dataIn[2410]),
.io_parallelIn_2411(dataIn[2411]),
.io_parallelIn_2412(dataIn[2412]),
.io_parallelIn_2413(dataIn[2413]),
.io_parallelIn_2414(dataIn[2414]),
.io_parallelIn_2415(dataIn[2415]),
.io_parallelIn_2416(dataIn[2416]),
.io_parallelIn_2417(dataIn[2417]),
.io_parallelIn_2418(dataIn[2418]),
.io_parallelIn_2419(dataIn[2419]),
.io_parallelIn_2420(dataIn[2420]),
.io_parallelIn_2421(dataIn[2421]),
.io_parallelIn_2422(dataIn[2422]),
.io_parallelIn_2423(dataIn[2423]),
.io_parallelIn_2424(dataIn[2424]),
.io_parallelIn_2425(dataIn[2425]),
.io_parallelIn_2426(dataIn[2426]),
.io_parallelIn_2427(dataIn[2427]),
.io_parallelIn_2428(dataIn[2428]),
.io_parallelIn_2429(dataIn[2429]),
.io_parallelIn_2430(dataIn[2430]),
.io_parallelIn_2431(dataIn[2431]),
.io_parallelIn_2432(dataIn[2432]),
.io_parallelIn_2433(dataIn[2433]),
.io_parallelIn_2434(dataIn[2434]),
.io_parallelIn_2435(dataIn[2435]),
.io_parallelIn_2436(dataIn[2436]),
.io_parallelIn_2437(dataIn[2437]),
.io_parallelIn_2438(dataIn[2438]),
.io_parallelIn_2439(dataIn[2439]),
.io_parallelIn_2440(dataIn[2440]),
.io_parallelIn_2441(dataIn[2441]),
.io_parallelIn_2442(dataIn[2442]),
.io_parallelIn_2443(dataIn[2443]),
.io_parallelIn_2444(dataIn[2444]),
.io_parallelIn_2445(dataIn[2445]),
.io_parallelIn_2446(dataIn[2446]),
.io_parallelIn_2447(dataIn[2447]),
.io_parallelIn_2448(dataIn[2448]),
.io_parallelIn_2449(dataIn[2449]),
.io_parallelIn_2450(dataIn[2450]),
.io_parallelIn_2451(dataIn[2451]),
.io_parallelIn_2452(dataIn[2452]),
.io_parallelIn_2453(dataIn[2453]),
.io_parallelIn_2454(dataIn[2454]),
.io_parallelIn_2455(dataIn[2455]),
.io_parallelIn_2456(dataIn[2456]),
.io_parallelIn_2457(dataIn[2457]),
.io_parallelIn_2458(dataIn[2458]),
.io_parallelIn_2459(dataIn[2459]),
.io_parallelIn_2460(dataIn[2460]),
.io_parallelIn_2461(dataIn[2461]),
.io_parallelIn_2462(dataIn[2462]),
.io_parallelIn_2463(dataIn[2463]),
.io_parallelIn_2464(dataIn[2464]),
.io_parallelIn_2465(dataIn[2465]),
.io_parallelIn_2466(dataIn[2466]),
.io_parallelIn_2467(dataIn[2467]),
.io_parallelIn_2468(dataIn[2468]),
.io_parallelIn_2469(dataIn[2469]),
.io_parallelIn_2470(dataIn[2470]),
.io_parallelIn_2471(dataIn[2471]),
.io_parallelIn_2472(dataIn[2472]),
.io_parallelIn_2473(dataIn[2473]),
.io_parallelIn_2474(dataIn[2474]),
.io_parallelIn_2475(dataIn[2475]),
.io_parallelIn_2476(dataIn[2476]),
.io_parallelIn_2477(dataIn[2477]),
.io_parallelIn_2478(dataIn[2478]),
.io_parallelIn_2479(dataIn[2479]),
.io_parallelIn_2480(dataIn[2480]),
.io_parallelIn_2481(dataIn[2481]),
.io_parallelIn_2482(dataIn[2482]),
.io_parallelIn_2483(dataIn[2483]),
.io_parallelIn_2484(dataIn[2484]),
.io_parallelIn_2485(dataIn[2485]),
.io_parallelIn_2486(dataIn[2486]),
.io_parallelIn_2487(dataIn[2487]),
.io_parallelIn_2488(dataIn[2488]),
.io_parallelIn_2489(dataIn[2489]),
.io_parallelIn_2490(dataIn[2490]),
.io_parallelIn_2491(dataIn[2491]),
.io_parallelIn_2492(dataIn[2492]),
.io_parallelIn_2493(dataIn[2493]),
.io_parallelIn_2494(dataIn[2494]),
.io_parallelIn_2495(dataIn[2495]),
.io_parallelIn_2496(dataIn[2496]),
.io_parallelIn_2497(dataIn[2497]),
.io_parallelIn_2498(dataIn[2498]),
.io_parallelIn_2499(dataIn[2499]),
.io_parallelIn_2500(dataIn[2500]),
.io_parallelIn_2501(dataIn[2501]),
.io_parallelIn_2502(dataIn[2502]),
.io_parallelIn_2503(dataIn[2503]),
.io_parallelIn_2504(dataIn[2504]),
.io_parallelIn_2505(dataIn[2505]),
.io_parallelIn_2506(dataIn[2506]),
.io_parallelIn_2507(dataIn[2507]),
.io_parallelIn_2508(dataIn[2508]),
.io_parallelIn_2509(dataIn[2509]),
.io_parallelIn_2510(dataIn[2510]),
.io_parallelIn_2511(dataIn[2511]),
.io_parallelIn_2512(dataIn[2512]),
.io_parallelIn_2513(dataIn[2513]),
.io_parallelIn_2514(dataIn[2514]),
.io_parallelIn_2515(dataIn[2515]),
.io_parallelIn_2516(dataIn[2516]),
.io_parallelIn_2517(dataIn[2517]),
.io_parallelIn_2518(dataIn[2518]),
.io_parallelIn_2519(dataIn[2519]),
.io_parallelIn_2520(dataIn[2520]),
.io_parallelIn_2521(dataIn[2521]),
.io_parallelIn_2522(dataIn[2522]),
.io_parallelIn_2523(dataIn[2523]),
.io_parallelIn_2524(dataIn[2524]),
.io_parallelIn_2525(dataIn[2525]),
.io_parallelIn_2526(dataIn[2526]),
.io_parallelIn_2527(dataIn[2527]),
.io_parallelIn_2528(dataIn[2528]),
.io_parallelIn_2529(dataIn[2529]),
.io_parallelIn_2530(dataIn[2530]),
.io_parallelIn_2531(dataIn[2531]),
.io_parallelIn_2532(dataIn[2532]),
.io_parallelIn_2533(dataIn[2533]),
.io_parallelIn_2534(dataIn[2534]),
.io_parallelIn_2535(dataIn[2535]),
.io_parallelIn_2536(dataIn[2536]),
.io_parallelIn_2537(dataIn[2537]),
.io_parallelIn_2538(dataIn[2538]),
.io_parallelIn_2539(dataIn[2539]),
.io_parallelIn_2540(dataIn[2540]),
.io_parallelIn_2541(dataIn[2541]),
.io_parallelIn_2542(dataIn[2542]),
.io_parallelIn_2543(dataIn[2543]),
.io_parallelIn_2544(dataIn[2544]),
.io_parallelIn_2545(dataIn[2545]),
.io_parallelIn_2546(dataIn[2546]),
.io_parallelIn_2547(dataIn[2547]),
.io_parallelIn_2548(dataIn[2548]),
.io_parallelIn_2549(dataIn[2549]),
.io_parallelIn_2550(dataIn[2550]),
.io_parallelIn_2551(dataIn[2551]),
.io_parallelIn_2552(dataIn[2552]),
.io_parallelIn_2553(dataIn[2553]),
.io_parallelIn_2554(dataIn[2554]),
.io_parallelIn_2555(dataIn[2555]),
.io_parallelIn_2556(dataIn[2556]),
.io_parallelIn_2557(dataIn[2557]),
.io_parallelIn_2558(dataIn[2558]),
.io_parallelIn_2559(dataIn[2559]),
.io_parallelIn_2560(dataIn[2560]),
.io_parallelIn_2561(dataIn[2561]),
.io_parallelIn_2562(dataIn[2562]),
.io_parallelIn_2563(dataIn[2563]),
.io_parallelIn_2564(dataIn[2564]),
.io_parallelIn_2565(dataIn[2565]),
.io_parallelIn_2566(dataIn[2566]),
.io_parallelIn_2567(dataIn[2567]),
.io_parallelIn_2568(dataIn[2568]),
.io_parallelIn_2569(dataIn[2569]),
.io_parallelIn_2570(dataIn[2570]),
.io_parallelIn_2571(dataIn[2571]),
.io_parallelIn_2572(dataIn[2572]),
.io_parallelIn_2573(dataIn[2573]),
.io_parallelIn_2574(dataIn[2574]),
.io_parallelIn_2575(dataIn[2575]),
.io_parallelIn_2576(dataIn[2576]),
.io_parallelIn_2577(dataIn[2577]),
.io_parallelIn_2578(dataIn[2578]),
.io_parallelIn_2579(dataIn[2579]),
.io_parallelIn_2580(dataIn[2580]),
.io_parallelIn_2581(dataIn[2581]),
.io_parallelIn_2582(dataIn[2582]),
.io_parallelIn_2583(dataIn[2583]),
.io_parallelIn_2584(dataIn[2584]),
.io_parallelIn_2585(dataIn[2585]),
.io_parallelIn_2586(dataIn[2586]),
.io_parallelIn_2587(dataIn[2587]),
.io_parallelIn_2588(dataIn[2588]),
.io_parallelIn_2589(dataIn[2589]),
.io_parallelIn_2590(dataIn[2590]),
.io_parallelIn_2591(dataIn[2591]),
.io_parallelIn_2592(dataIn[2592]),
.io_parallelIn_2593(dataIn[2593]),
.io_parallelIn_2594(dataIn[2594]),
.io_parallelIn_2595(dataIn[2595]),
.io_parallelIn_2596(dataIn[2596]),
.io_parallelIn_2597(dataIn[2597]),
.io_parallelIn_2598(dataIn[2598]),
.io_parallelIn_2599(dataIn[2599]),
.io_parallelIn_2600(dataIn[2600]),
.io_parallelIn_2601(dataIn[2601]),
.io_parallelIn_2602(dataIn[2602]),
.io_parallelIn_2603(dataIn[2603]),
.io_parallelIn_2604(dataIn[2604]),
.io_parallelIn_2605(dataIn[2605]),
.io_parallelIn_2606(dataIn[2606]),
.io_parallelIn_2607(dataIn[2607]),
.io_parallelIn_2608(dataIn[2608]),
.io_parallelIn_2609(dataIn[2609]),
.io_parallelIn_2610(dataIn[2610]),
.io_parallelIn_2611(dataIn[2611]),
.io_parallelIn_2612(dataIn[2612]),
.io_parallelIn_2613(dataIn[2613]),
.io_parallelIn_2614(dataIn[2614]),
.io_parallelIn_2615(dataIn[2615]),
.io_parallelIn_2616(dataIn[2616]),
.io_parallelIn_2617(dataIn[2617]),
.io_parallelIn_2618(dataIn[2618]),
.io_parallelIn_2619(dataIn[2619]),
.io_parallelIn_2620(dataIn[2620]),
.io_parallelIn_2621(dataIn[2621]),
.io_parallelIn_2622(dataIn[2622]),
.io_parallelIn_2623(dataIn[2623]),
.io_parallelIn_2624(dataIn[2624]),
.io_parallelIn_2625(dataIn[2625]),
.io_parallelIn_2626(dataIn[2626]),
.io_parallelIn_2627(dataIn[2627]),
.io_parallelIn_2628(dataIn[2628]),
.io_parallelIn_2629(dataIn[2629]),
.io_parallelIn_2630(dataIn[2630]),
.io_parallelIn_2631(dataIn[2631]),
.io_parallelIn_2632(dataIn[2632]),
.io_parallelIn_2633(dataIn[2633]),
.io_parallelIn_2634(dataIn[2634]),
.io_parallelIn_2635(dataIn[2635]),
.io_parallelIn_2636(dataIn[2636]),
.io_parallelIn_2637(dataIn[2637]),
.io_parallelIn_2638(dataIn[2638]),
.io_parallelIn_2639(dataIn[2639]),
.io_parallelIn_2640(dataIn[2640]),
.io_parallelIn_2641(dataIn[2641]),
.io_parallelIn_2642(dataIn[2642]),
.io_parallelIn_2643(dataIn[2643]),
.io_parallelIn_2644(dataIn[2644]),
.io_parallelIn_2645(dataIn[2645]),
.io_parallelIn_2646(dataIn[2646]),
.io_parallelIn_2647(dataIn[2647]),
.io_parallelIn_2648(dataIn[2648]),
.io_parallelIn_2649(dataIn[2649]),
.io_parallelIn_2650(dataIn[2650]),
.io_parallelIn_2651(dataIn[2651]),
.io_parallelIn_2652(dataIn[2652]),
.io_parallelIn_2653(dataIn[2653]),
.io_parallelIn_2654(dataIn[2654]),
.io_parallelIn_2655(dataIn[2655]),
.io_parallelIn_2656(dataIn[2656]),
.io_parallelIn_2657(dataIn[2657]),
.io_parallelIn_2658(dataIn[2658]),
.io_parallelIn_2659(dataIn[2659]),
.io_parallelIn_2660(dataIn[2660]),
.io_parallelIn_2661(dataIn[2661]),
.io_parallelIn_2662(dataIn[2662]),
.io_parallelIn_2663(dataIn[2663]),
.io_parallelIn_2664(dataIn[2664]),
.io_parallelIn_2665(dataIn[2665]),
.io_parallelIn_2666(dataIn[2666]),
.io_parallelIn_2667(dataIn[2667]),
.io_parallelIn_2668(dataIn[2668]),
.io_parallelIn_2669(dataIn[2669]),
.io_parallelIn_2670(dataIn[2670]),
.io_parallelIn_2671(dataIn[2671]),
.io_parallelIn_2672(dataIn[2672]),
.io_parallelIn_2673(dataIn[2673]),
.io_parallelIn_2674(dataIn[2674]),
.io_parallelIn_2675(dataIn[2675]),
.io_parallelIn_2676(dataIn[2676]),
.io_parallelIn_2677(dataIn[2677]),
.io_parallelIn_2678(dataIn[2678]),
.io_parallelIn_2679(dataIn[2679]),
.io_parallelIn_2680(dataIn[2680]),
.io_parallelIn_2681(dataIn[2681]),
.io_parallelIn_2682(dataIn[2682]),
.io_parallelIn_2683(dataIn[2683]),
.io_parallelIn_2684(dataIn[2684]),
.io_parallelIn_2685(dataIn[2685]),
.io_parallelIn_2686(dataIn[2686]),
.io_parallelIn_2687(dataIn[2687]),
.io_parallelIn_2688(dataIn[2688]),
.io_parallelIn_2689(dataIn[2689]),
.io_parallelIn_2690(dataIn[2690]),
.io_parallelIn_2691(dataIn[2691]),
.io_parallelIn_2692(dataIn[2692]),
.io_parallelIn_2693(dataIn[2693]),
.io_parallelIn_2694(dataIn[2694]),
.io_parallelIn_2695(dataIn[2695]),
.io_parallelIn_2696(dataIn[2696]),
.io_parallelIn_2697(dataIn[2697]),
.io_parallelIn_2698(dataIn[2698]),
.io_parallelIn_2699(dataIn[2699]),
.io_parallelIn_2700(dataIn[2700]),
.io_parallelIn_2701(dataIn[2701]),
.io_parallelIn_2702(dataIn[2702]),
.io_parallelIn_2703(dataIn[2703]),
.io_parallelIn_2704(dataIn[2704]),
.io_parallelIn_2705(dataIn[2705]),
.io_parallelIn_2706(dataIn[2706]),
.io_parallelIn_2707(dataIn[2707]),
.io_parallelIn_2708(dataIn[2708]),
.io_parallelIn_2709(dataIn[2709]),
.io_parallelIn_2710(dataIn[2710]),
.io_parallelIn_2711(dataIn[2711]),
.io_parallelIn_2712(dataIn[2712]),
.io_parallelIn_2713(dataIn[2713]),
.io_parallelIn_2714(dataIn[2714]),
.io_parallelIn_2715(dataIn[2715]),
.io_parallelIn_2716(dataIn[2716]),
.io_parallelIn_2717(dataIn[2717]),
.io_parallelIn_2718(dataIn[2718]),
.io_parallelIn_2719(dataIn[2719]),
.io_parallelIn_2720(dataIn[2720]),
.io_parallelIn_2721(dataIn[2721]),
.io_parallelIn_2722(dataIn[2722]),
.io_parallelIn_2723(dataIn[2723]),
.io_parallelIn_2724(dataIn[2724]),
.io_parallelIn_2725(dataIn[2725]),
.io_parallelIn_2726(dataIn[2726]),
.io_parallelIn_2727(dataIn[2727]),
.io_parallelIn_2728(dataIn[2728]),
.io_parallelIn_2729(dataIn[2729]),
.io_parallelIn_2730(dataIn[2730]),
.io_parallelIn_2731(dataIn[2731]),
.io_parallelIn_2732(dataIn[2732]),
.io_parallelIn_2733(dataIn[2733]),
.io_parallelIn_2734(dataIn[2734]),
.io_parallelIn_2735(dataIn[2735]),
.io_parallelIn_2736(dataIn[2736]),
.io_parallelIn_2737(dataIn[2737]),
.io_parallelIn_2738(dataIn[2738]),
.io_parallelIn_2739(dataIn[2739]),
.io_parallelIn_2740(dataIn[2740]),
.io_parallelIn_2741(dataIn[2741]),
.io_parallelIn_2742(dataIn[2742]),
.io_parallelIn_2743(dataIn[2743]),
.io_parallelIn_2744(dataIn[2744]),
.io_parallelIn_2745(dataIn[2745]),
.io_parallelIn_2746(dataIn[2746]),
.io_parallelIn_2747(dataIn[2747]),
.io_parallelIn_2748(dataIn[2748]),
.io_parallelIn_2749(dataIn[2749]),
.io_parallelIn_2750(dataIn[2750]),
.io_parallelIn_2751(dataIn[2751]),
.io_parallelIn_2752(dataIn[2752]),
.io_parallelIn_2753(dataIn[2753]),
.io_parallelIn_2754(dataIn[2754]),
.io_parallelIn_2755(dataIn[2755]),
.io_parallelIn_2756(dataIn[2756]),
.io_parallelIn_2757(dataIn[2757]),
.io_parallelIn_2758(dataIn[2758]),
.io_parallelIn_2759(dataIn[2759]),
.io_parallelIn_2760(dataIn[2760]),
.io_parallelIn_2761(dataIn[2761]),
.io_parallelIn_2762(dataIn[2762]),
.io_parallelIn_2763(dataIn[2763]),
.io_parallelIn_2764(dataIn[2764]),
.io_parallelIn_2765(dataIn[2765]),
.io_parallelIn_2766(dataIn[2766]),
.io_parallelIn_2767(dataIn[2767]),
.io_parallelIn_2768(dataIn[2768]),
.io_parallelIn_2769(dataIn[2769]),
.io_parallelIn_2770(dataIn[2770]),
.io_parallelIn_2771(dataIn[2771]),
.io_parallelIn_2772(dataIn[2772]),
.io_parallelIn_2773(dataIn[2773]),
.io_parallelIn_2774(dataIn[2774]),
.io_parallelIn_2775(dataIn[2775]),
.io_parallelIn_2776(dataIn[2776]),
.io_parallelIn_2777(dataIn[2777]),
.io_parallelIn_2778(dataIn[2778]),
.io_parallelIn_2779(dataIn[2779]),
.io_parallelIn_2780(dataIn[2780]),
.io_parallelIn_2781(dataIn[2781]),
.io_parallelIn_2782(dataIn[2782]),
.io_parallelIn_2783(dataIn[2783]),
.io_parallelIn_2784(dataIn[2784]),
.io_parallelIn_2785(dataIn[2785]),
.io_parallelIn_2786(dataIn[2786]),
.io_parallelIn_2787(dataIn[2787]),
.io_parallelIn_2788(dataIn[2788]),
.io_parallelIn_2789(dataIn[2789]),
.io_parallelIn_2790(dataIn[2790]),
.io_parallelIn_2791(dataIn[2791]),
.io_parallelIn_2792(dataIn[2792]),
.io_parallelIn_2793(dataIn[2793]),
.io_parallelIn_2794(dataIn[2794]),
.io_parallelIn_2795(dataIn[2795]),
.io_parallelIn_2796(dataIn[2796]),
.io_parallelIn_2797(dataIn[2797]),
.io_parallelIn_2798(dataIn[2798]),
.io_parallelIn_2799(dataIn[2799]),
.io_parallelIn_2800(dataIn[2800]),
.io_parallelIn_2801(dataIn[2801]),
.io_parallelIn_2802(dataIn[2802]),
.io_parallelIn_2803(dataIn[2803]),
.io_parallelIn_2804(dataIn[2804]),
.io_parallelIn_2805(dataIn[2805]),
.io_parallelIn_2806(dataIn[2806]),
.io_parallelIn_2807(dataIn[2807]),
.io_parallelIn_2808(dataIn[2808]),
.io_parallelIn_2809(dataIn[2809]),
.io_parallelIn_2810(dataIn[2810]),
.io_parallelIn_2811(dataIn[2811]),
.io_parallelIn_2812(dataIn[2812]),
.io_parallelIn_2813(dataIn[2813]),
.io_parallelIn_2814(dataIn[2814]),
.io_parallelIn_2815(dataIn[2815]),
.io_parallelIn_2816(dataIn[2816]),
.io_parallelIn_2817(dataIn[2817]),
.io_parallelIn_2818(dataIn[2818]),
.io_parallelIn_2819(dataIn[2819]),
.io_parallelIn_2820(dataIn[2820]),
.io_parallelIn_2821(dataIn[2821]),
.io_parallelIn_2822(dataIn[2822]),
.io_parallelIn_2823(dataIn[2823]),
.io_parallelIn_2824(dataIn[2824]),
.io_parallelIn_2825(dataIn[2825]),
.io_parallelIn_2826(dataIn[2826]),
.io_parallelIn_2827(dataIn[2827]),
.io_parallelIn_2828(dataIn[2828]),
.io_parallelIn_2829(dataIn[2829]),
.io_parallelIn_2830(dataIn[2830]),
.io_parallelIn_2831(dataIn[2831]),
.io_parallelIn_2832(dataIn[2832]),
.io_parallelIn_2833(dataIn[2833]),
.io_parallelIn_2834(dataIn[2834]),
.io_parallelIn_2835(dataIn[2835]),
.io_parallelIn_2836(dataIn[2836]),
.io_parallelIn_2837(dataIn[2837]),
.io_parallelIn_2838(dataIn[2838]),
.io_parallelIn_2839(dataIn[2839]),
.io_parallelIn_2840(dataIn[2840]),
.io_parallelIn_2841(dataIn[2841]),
.io_parallelIn_2842(dataIn[2842]),
.io_parallelIn_2843(dataIn[2843]),
.io_parallelIn_2844(dataIn[2844]),
.io_parallelIn_2845(dataIn[2845]),
.io_parallelIn_2846(dataIn[2846]),
.io_parallelIn_2847(dataIn[2847]),
.io_parallelIn_2848(dataIn[2848]),
.io_parallelIn_2849(dataIn[2849]),
.io_parallelIn_2850(dataIn[2850]),
.io_parallelIn_2851(dataIn[2851]),
.io_parallelIn_2852(dataIn[2852]),
.io_parallelIn_2853(dataIn[2853]),
.io_parallelIn_2854(dataIn[2854]),
.io_parallelIn_2855(dataIn[2855]),
.io_parallelIn_2856(dataIn[2856]),
.io_parallelIn_2857(dataIn[2857]),
.io_parallelIn_2858(dataIn[2858]),
.io_parallelIn_2859(dataIn[2859]),
.io_parallelIn_2860(dataIn[2860]),
.io_parallelIn_2861(dataIn[2861]),
.io_parallelIn_2862(dataIn[2862]),
.io_parallelIn_2863(dataIn[2863]),
.io_parallelIn_2864(dataIn[2864]),
.io_parallelIn_2865(dataIn[2865]),
.io_parallelIn_2866(dataIn[2866]),
.io_parallelIn_2867(dataIn[2867]),
.io_parallelIn_2868(dataIn[2868]),
.io_parallelIn_2869(dataIn[2869]),
.io_parallelIn_2870(dataIn[2870]),
.io_parallelIn_2871(dataIn[2871]),
.io_parallelIn_2872(dataIn[2872]),
.io_parallelIn_2873(dataIn[2873]),
.io_parallelIn_2874(dataIn[2874]),
.io_parallelIn_2875(dataIn[2875]),
.io_parallelIn_2876(dataIn[2876]),
.io_parallelIn_2877(dataIn[2877]),
.io_parallelIn_2878(dataIn[2878]),
.io_parallelIn_2879(dataIn[2879]),
.io_parallelIn_2880(dataIn[2880]),
.io_parallelIn_2881(dataIn[2881]),
.io_parallelIn_2882(dataIn[2882]),
.io_parallelIn_2883(dataIn[2883]),
.io_parallelIn_2884(dataIn[2884]),
.io_parallelIn_2885(dataIn[2885]),
.io_parallelIn_2886(dataIn[2886]),
.io_parallelIn_2887(dataIn[2887]),
.io_parallelIn_2888(dataIn[2888]),
.io_parallelIn_2889(dataIn[2889]),
.io_parallelIn_2890(dataIn[2890]),
.io_parallelIn_2891(dataIn[2891]),
.io_parallelIn_2892(dataIn[2892]),
.io_parallelIn_2893(dataIn[2893]),
.io_parallelIn_2894(dataIn[2894]),
.io_parallelIn_2895(dataIn[2895]),
.io_parallelIn_2896(dataIn[2896]),
.io_parallelIn_2897(dataIn[2897]),
.io_parallelIn_2898(dataIn[2898]),
.io_parallelIn_2899(dataIn[2899]),
.io_parallelIn_2900(dataIn[2900]),
.io_parallelIn_2901(dataIn[2901]),
.io_parallelIn_2902(dataIn[2902]),
.io_parallelIn_2903(dataIn[2903]),
.io_parallelIn_2904(dataIn[2904]),
.io_parallelIn_2905(dataIn[2905]),
.io_parallelIn_2906(dataIn[2906]),
.io_parallelIn_2907(dataIn[2907]),
.io_parallelIn_2908(dataIn[2908]),
.io_parallelIn_2909(dataIn[2909]),
.io_parallelIn_2910(dataIn[2910]),
.io_parallelIn_2911(dataIn[2911]),
.io_parallelIn_2912(dataIn[2912]),
.io_parallelIn_2913(dataIn[2913]),
.io_parallelIn_2914(dataIn[2914]),
.io_parallelIn_2915(dataIn[2915]),
.io_parallelIn_2916(dataIn[2916]),
.io_parallelIn_2917(dataIn[2917]),
.io_parallelIn_2918(dataIn[2918]),
.io_parallelIn_2919(dataIn[2919]),
.io_parallelIn_2920(dataIn[2920]),
.io_parallelIn_2921(dataIn[2921]),
.io_parallelIn_2922(dataIn[2922]),
.io_parallelIn_2923(dataIn[2923]),
.io_parallelIn_2924(dataIn[2924]),
.io_parallelIn_2925(dataIn[2925]),
.io_parallelIn_2926(dataIn[2926]),
.io_parallelIn_2927(dataIn[2927]),
.io_parallelIn_2928(dataIn[2928]),
.io_parallelIn_2929(dataIn[2929]),
.io_parallelIn_2930(dataIn[2930]),
.io_parallelIn_2931(dataIn[2931]),
.io_parallelIn_2932(dataIn[2932]),
.io_parallelIn_2933(dataIn[2933]),
.io_parallelIn_2934(dataIn[2934]),
.io_parallelIn_2935(dataIn[2935]),
.io_parallelIn_2936(dataIn[2936]),
.io_parallelIn_2937(dataIn[2937]),
.io_parallelIn_2938(dataIn[2938]),
.io_parallelIn_2939(dataIn[2939]),
.io_parallelIn_2940(dataIn[2940]),
.io_parallelIn_2941(dataIn[2941]),
.io_parallelIn_2942(dataIn[2942]),
.io_parallelIn_2943(dataIn[2943]),
.io_parallelIn_2944(dataIn[2944]),
.io_parallelIn_2945(dataIn[2945]),
.io_parallelIn_2946(dataIn[2946]),
.io_parallelIn_2947(dataIn[2947]),
.io_parallelIn_2948(dataIn[2948]),
.io_parallelIn_2949(dataIn[2949]),
.io_parallelIn_2950(dataIn[2950]),
.io_parallelIn_2951(dataIn[2951]),
.io_parallelIn_2952(dataIn[2952]),
.io_parallelIn_2953(dataIn[2953]),
.io_parallelIn_2954(dataIn[2954]),
.io_parallelIn_2955(dataIn[2955]),
.io_parallelIn_2956(dataIn[2956]),
.io_parallelIn_2957(dataIn[2957]),
.io_parallelIn_2958(dataIn[2958]),
.io_parallelIn_2959(dataIn[2959]),
.io_parallelIn_2960(dataIn[2960]),
.io_parallelIn_2961(dataIn[2961]),
.io_parallelIn_2962(dataIn[2962]),
.io_parallelIn_2963(dataIn[2963]),
.io_parallelIn_2964(dataIn[2964]),
.io_parallelIn_2965(dataIn[2965]),
.io_parallelIn_2966(dataIn[2966]),
.io_parallelIn_2967(dataIn[2967]),
.io_parallelIn_2968(dataIn[2968]),
.io_parallelIn_2969(dataIn[2969]),
.io_parallelIn_2970(dataIn[2970]),
.io_parallelIn_2971(dataIn[2971]),
.io_parallelIn_2972(dataIn[2972]),
.io_parallelIn_2973(dataIn[2973]),
.io_parallelIn_2974(dataIn[2974]),
.io_parallelIn_2975(dataIn[2975]),
.io_parallelIn_2976(dataIn[2976]),
.io_parallelIn_2977(dataIn[2977]),
.io_parallelIn_2978(dataIn[2978]),
.io_parallelIn_2979(dataIn[2979]),
.io_parallelIn_2980(dataIn[2980]),
.io_parallelIn_2981(dataIn[2981]),
.io_parallelIn_2982(dataIn[2982]),
.io_parallelIn_2983(dataIn[2983]),
.io_parallelIn_2984(dataIn[2984]),
.io_parallelIn_2985(dataIn[2985]),
.io_parallelIn_2986(dataIn[2986]),
.io_parallelIn_2987(dataIn[2987]),
.io_parallelIn_2988(dataIn[2988]),
.io_parallelIn_2989(dataIn[2989]),
.io_parallelIn_2990(dataIn[2990]),
.io_parallelIn_2991(dataIn[2991]),
.io_parallelIn_2992(dataIn[2992]),
.io_parallelIn_2993(dataIn[2993]),
.io_parallelIn_2994(dataIn[2994]),
.io_parallelIn_2995(dataIn[2995]),
.io_parallelIn_2996(dataIn[2996]),
.io_parallelIn_2997(dataIn[2997]),
.io_parallelIn_2998(dataIn[2998]),
.io_parallelIn_2999(dataIn[2999]),
.io_parallelIn_3000(dataIn[3000]),
.io_parallelIn_3001(dataIn[3001]),
.io_parallelIn_3002(dataIn[3002]),
.io_parallelIn_3003(dataIn[3003]),
.io_parallelIn_3004(dataIn[3004]),
.io_parallelIn_3005(dataIn[3005]),
.io_parallelIn_3006(dataIn[3006]),
.io_parallelIn_3007(dataIn[3007]),
.io_parallelIn_3008(dataIn[3008]),
.io_parallelIn_3009(dataIn[3009]),
.io_parallelIn_3010(dataIn[3010]),
.io_parallelIn_3011(dataIn[3011]),
.io_parallelIn_3012(dataIn[3012]),
.io_parallelIn_3013(dataIn[3013]),
.io_parallelIn_3014(dataIn[3014]),
.io_parallelIn_3015(dataIn[3015]),
.io_parallelIn_3016(dataIn[3016]),
.io_parallelIn_3017(dataIn[3017]),
.io_parallelIn_3018(dataIn[3018]),
.io_parallelIn_3019(dataIn[3019]),
.io_parallelIn_3020(dataIn[3020]),
.io_parallelIn_3021(dataIn[3021]),
.io_parallelIn_3022(dataIn[3022]),
.io_parallelIn_3023(dataIn[3023]),
.io_parallelIn_3024(dataIn[3024]),
.io_parallelIn_3025(dataIn[3025]),
.io_parallelIn_3026(dataIn[3026]),
.io_parallelIn_3027(dataIn[3027]),
.io_parallelIn_3028(dataIn[3028]),
.io_parallelIn_3029(dataIn[3029]),
.io_parallelIn_3030(dataIn[3030]),
.io_parallelIn_3031(dataIn[3031]),
.io_parallelIn_3032(dataIn[3032]),
.io_parallelIn_3033(dataIn[3033]),
.io_parallelIn_3034(dataIn[3034]),
.io_parallelIn_3035(dataIn[3035]),
.io_parallelIn_3036(dataIn[3036]),
.io_parallelIn_3037(dataIn[3037]),
.io_parallelIn_3038(dataIn[3038]),
.io_parallelIn_3039(dataIn[3039]),
.io_parallelIn_3040(dataIn[3040]),
.io_parallelIn_3041(dataIn[3041]),
.io_parallelIn_3042(dataIn[3042]),
.io_parallelIn_3043(dataIn[3043]),
.io_parallelIn_3044(dataIn[3044]),
.io_parallelIn_3045(dataIn[3045]),
.io_parallelIn_3046(dataIn[3046]),
.io_parallelIn_3047(dataIn[3047]),
.io_parallelIn_3048(dataIn[3048]),
.io_parallelIn_3049(dataIn[3049]),
.io_parallelIn_3050(dataIn[3050]),
.io_parallelIn_3051(dataIn[3051]),
.io_parallelIn_3052(dataIn[3052]),
.io_parallelIn_3053(dataIn[3053]),
.io_parallelIn_3054(dataIn[3054]),
.io_parallelIn_3055(dataIn[3055]),
.io_parallelIn_3056(dataIn[3056]),
.io_parallelIn_3057(dataIn[3057]),
.io_parallelIn_3058(dataIn[3058]),
.io_parallelIn_3059(dataIn[3059]),
.io_parallelIn_3060(dataIn[3060]),
.io_parallelIn_3061(dataIn[3061]),
.io_parallelIn_3062(dataIn[3062]),
.io_parallelIn_3063(dataIn[3063]),
.io_parallelIn_3064(dataIn[3064]),
.io_parallelIn_3065(dataIn[3065]),
.io_parallelIn_3066(dataIn[3066]),
.io_parallelIn_3067(dataIn[3067]),
.io_parallelIn_3068(dataIn[3068]),
.io_parallelIn_3069(dataIn[3069]),
.io_parallelIn_3070(dataIn[3070]),
.io_parallelIn_3071(dataIn[3071]),
.io_parallelIn_3072(dataIn[3072]),
.io_parallelIn_3073(dataIn[3073]),
.io_parallelIn_3074(dataIn[3074]),
.io_parallelIn_3075(dataIn[3075]),
.io_parallelIn_3076(dataIn[3076]),
.io_parallelIn_3077(dataIn[3077]),
.io_parallelIn_3078(dataIn[3078]),
.io_parallelIn_3079(dataIn[3079]),
.io_parallelIn_3080(dataIn[3080]),
.io_parallelIn_3081(dataIn[3081]),
.io_parallelIn_3082(dataIn[3082]),
.io_parallelIn_3083(dataIn[3083]),
.io_parallelIn_3084(dataIn[3084]),
.io_parallelIn_3085(dataIn[3085]),
.io_parallelIn_3086(dataIn[3086]),
.io_parallelIn_3087(dataIn[3087]),
.io_parallelIn_3088(dataIn[3088]),
.io_parallelIn_3089(dataIn[3089]),
.io_parallelIn_3090(dataIn[3090]),
.io_parallelIn_3091(dataIn[3091]),
.io_parallelIn_3092(dataIn[3092]),
.io_parallelIn_3093(dataIn[3093]),
.io_parallelIn_3094(dataIn[3094]),
.io_parallelIn_3095(dataIn[3095]),
.io_parallelIn_3096(dataIn[3096]),
.io_parallelIn_3097(dataIn[3097]),
.io_parallelIn_3098(dataIn[3098]),
.io_parallelIn_3099(dataIn[3099]),
.io_parallelIn_3100(dataIn[3100]),
.io_parallelIn_3101(dataIn[3101]),
.io_parallelIn_3102(dataIn[3102]),
.io_parallelIn_3103(dataIn[3103]),
.io_parallelIn_3104(dataIn[3104]),
.io_parallelIn_3105(dataIn[3105]),
.io_parallelIn_3106(dataIn[3106]),
.io_parallelIn_3107(dataIn[3107]),
.io_parallelIn_3108(dataIn[3108]),
.io_parallelIn_3109(dataIn[3109]),
.io_parallelIn_3110(dataIn[3110]),
.io_parallelIn_3111(dataIn[3111]),
.io_parallelIn_3112(dataIn[3112]),
.io_parallelIn_3113(dataIn[3113]),
.io_parallelIn_3114(dataIn[3114]),
.io_parallelIn_3115(dataIn[3115]),
.io_parallelIn_3116(dataIn[3116]),
.io_parallelIn_3117(dataIn[3117]),
.io_parallelIn_3118(dataIn[3118]),
.io_parallelIn_3119(dataIn[3119]),
.io_parallelIn_3120(dataIn[3120]),
.io_parallelIn_3121(dataIn[3121]),
.io_parallelIn_3122(dataIn[3122]),
.io_parallelIn_3123(dataIn[3123]),
.io_parallelIn_3124(dataIn[3124]),
.io_parallelIn_3125(dataIn[3125]),
.io_parallelIn_3126(dataIn[3126]),
.io_parallelIn_3127(dataIn[3127]),
.io_parallelIn_3128(dataIn[3128]),
.io_parallelIn_3129(dataIn[3129]),
.io_parallelIn_3130(dataIn[3130]),
.io_parallelIn_3131(dataIn[3131]),
.io_parallelIn_3132(dataIn[3132]),
.io_parallelIn_3133(dataIn[3133]),
.io_parallelIn_3134(dataIn[3134]),
.io_parallelIn_3135(dataIn[3135]),
.io_parallelIn_3136(dataIn[3136]),
.io_parallelIn_3137(dataIn[3137]),
.io_parallelIn_3138(dataIn[3138]),
.io_parallelIn_3139(dataIn[3139]),
.io_parallelIn_3140(dataIn[3140]),
.io_parallelIn_3141(dataIn[3141]),
.io_parallelIn_3142(dataIn[3142]),
.io_parallelIn_3143(dataIn[3143]),
.io_parallelIn_3144(dataIn[3144]),
.io_parallelIn_3145(dataIn[3145]),
.io_parallelIn_3146(dataIn[3146]),
.io_parallelIn_3147(dataIn[3147]),
.io_parallelIn_3148(dataIn[3148]),
.io_parallelIn_3149(dataIn[3149]),
.io_parallelIn_3150(dataIn[3150]),
.io_parallelIn_3151(dataIn[3151]),
.io_parallelIn_3152(dataIn[3152]),
.io_parallelIn_3153(dataIn[3153]),
.io_parallelIn_3154(dataIn[3154]),
.io_parallelIn_3155(dataIn[3155]),
.io_parallelIn_3156(dataIn[3156]),
.io_parallelIn_3157(dataIn[3157]),
.io_parallelIn_3158(dataIn[3158]),
.io_parallelIn_3159(dataIn[3159]),
.io_parallelIn_3160(dataIn[3160]),
.io_parallelIn_3161(dataIn[3161]),
.io_parallelIn_3162(dataIn[3162]),
.io_parallelIn_3163(dataIn[3163]),
.io_parallelIn_3164(dataIn[3164]),
.io_parallelIn_3165(dataIn[3165]),
.io_parallelIn_3166(dataIn[3166]),
.io_parallelIn_3167(dataIn[3167]),
.io_parallelIn_3168(dataIn[3168]),
.io_parallelIn_3169(dataIn[3169]),
.io_parallelIn_3170(dataIn[3170]),
.io_parallelIn_3171(dataIn[3171]),
.io_parallelIn_3172(dataIn[3172]),
.io_parallelIn_3173(dataIn[3173]),
.io_parallelIn_3174(dataIn[3174]),
.io_parallelIn_3175(dataIn[3175]),
.io_parallelIn_3176(dataIn[3176]),
.io_parallelIn_3177(dataIn[3177]),
.io_parallelIn_3178(dataIn[3178]),
.io_parallelIn_3179(dataIn[3179]),
.io_parallelIn_3180(dataIn[3180]),
.io_parallelIn_3181(dataIn[3181]),
.io_parallelIn_3182(dataIn[3182]),
.io_parallelIn_3183(dataIn[3183]),
.io_parallelIn_3184(dataIn[3184]),
.io_parallelIn_3185(dataIn[3185]),
.io_parallelIn_3186(dataIn[3186]),
.io_parallelIn_3187(dataIn[3187]),
.io_parallelIn_3188(dataIn[3188]),
.io_parallelIn_3189(dataIn[3189]),
.io_parallelIn_3190(dataIn[3190]),
.io_parallelIn_3191(dataIn[3191]),
.io_parallelIn_3192(dataIn[3192]),
.io_parallelIn_3193(dataIn[3193]),
.io_parallelIn_3194(dataIn[3194]),
.io_parallelIn_3195(dataIn[3195]),
.io_parallelIn_3196(dataIn[3196]),
.io_parallelIn_3197(dataIn[3197]),
.io_parallelIn_3198(dataIn[3198]),
.io_parallelIn_3199(dataIn[3199]),
.io_parallelIn_3200(dataIn[3200]),
.io_parallelIn_3201(dataIn[3201]),
.io_parallelIn_3202(dataIn[3202]),
.io_parallelIn_3203(dataIn[3203]),
.io_parallelIn_3204(dataIn[3204]),
.io_parallelIn_3205(dataIn[3205]),
.io_parallelIn_3206(dataIn[3206]),
.io_parallelIn_3207(dataIn[3207]),
.io_parallelIn_3208(dataIn[3208]),
.io_parallelIn_3209(dataIn[3209]),
.io_parallelIn_3210(dataIn[3210]),
.io_parallelIn_3211(dataIn[3211]),
.io_parallelIn_3212(dataIn[3212]),
.io_parallelIn_3213(dataIn[3213]),
.io_parallelIn_3214(dataIn[3214]),
.io_parallelIn_3215(dataIn[3215]),
.io_parallelIn_3216(dataIn[3216]),
.io_parallelIn_3217(dataIn[3217]),
.io_parallelIn_3218(dataIn[3218]),
.io_parallelIn_3219(dataIn[3219]),
.io_parallelIn_3220(dataIn[3220]),
.io_parallelIn_3221(dataIn[3221]),
.io_parallelIn_3222(dataIn[3222]),
.io_parallelIn_3223(dataIn[3223]),
.io_parallelIn_3224(dataIn[3224]),
.io_parallelIn_3225(dataIn[3225]),
.io_parallelIn_3226(dataIn[3226]),
.io_parallelIn_3227(dataIn[3227]),
.io_parallelIn_3228(dataIn[3228]),
.io_parallelIn_3229(dataIn[3229]),
.io_parallelIn_3230(dataIn[3230]),
.io_parallelIn_3231(dataIn[3231]),
.io_parallelIn_3232(dataIn[3232]),
.io_parallelIn_3233(dataIn[3233]),
.io_parallelIn_3234(dataIn[3234]),
.io_parallelIn_3235(dataIn[3235]),
.io_parallelIn_3236(dataIn[3236]),
.io_parallelIn_3237(dataIn[3237]),
.io_parallelIn_3238(dataIn[3238]),
.io_parallelIn_3239(dataIn[3239]),
.io_parallelIn_3240(dataIn[3240]),
.io_parallelIn_3241(dataIn[3241]),
.io_parallelIn_3242(dataIn[3242]),
.io_parallelIn_3243(dataIn[3243]),
.io_parallelIn_3244(dataIn[3244]),
.io_parallelIn_3245(dataIn[3245]),
.io_parallelIn_3246(dataIn[3246]),
.io_parallelIn_3247(dataIn[3247]),
.io_parallelIn_3248(dataIn[3248]),
.io_parallelIn_3249(dataIn[3249]),
.io_parallelIn_3250(dataIn[3250]),
.io_parallelIn_3251(dataIn[3251]),
.io_parallelIn_3252(dataIn[3252]),
.io_parallelIn_3253(dataIn[3253]),
.io_parallelIn_3254(dataIn[3254]),
.io_parallelIn_3255(dataIn[3255]),
.io_parallelIn_3256(dataIn[3256]),
.io_parallelIn_3257(dataIn[3257]),
.io_parallelIn_3258(dataIn[3258]),
.io_parallelIn_3259(dataIn[3259]),
.io_parallelIn_3260(dataIn[3260]),
.io_parallelIn_3261(dataIn[3261]),
.io_parallelIn_3262(dataIn[3262]),
.io_parallelIn_3263(dataIn[3263]),
.io_parallelIn_3264(dataIn[3264]),
.io_parallelIn_3265(dataIn[3265]),
.io_parallelIn_3266(dataIn[3266]),
.io_parallelIn_3267(dataIn[3267]),
.io_parallelIn_3268(dataIn[3268]),
.io_parallelIn_3269(dataIn[3269]),
.io_parallelIn_3270(dataIn[3270]),
.io_parallelIn_3271(dataIn[3271]),
.io_parallelIn_3272(dataIn[3272]),
.io_parallelIn_3273(dataIn[3273]),
.io_parallelIn_3274(dataIn[3274]),
.io_parallelIn_3275(dataIn[3275]),
.io_parallelIn_3276(dataIn[3276]),
.io_parallelIn_3277(dataIn[3277]),
.io_parallelIn_3278(dataIn[3278]),
.io_parallelIn_3279(dataIn[3279]),
.io_parallelIn_3280(dataIn[3280]),
.io_parallelIn_3281(dataIn[3281]),
.io_parallelIn_3282(dataIn[3282]),
.io_parallelIn_3283(dataIn[3283]),
.io_parallelIn_3284(dataIn[3284]),
.io_parallelIn_3285(dataIn[3285]),
.io_parallelIn_3286(dataIn[3286]),
.io_parallelIn_3287(dataIn[3287]),
.io_parallelIn_3288(dataIn[3288]),
.io_parallelIn_3289(dataIn[3289]),
.io_parallelIn_3290(dataIn[3290]),
.io_parallelIn_3291(dataIn[3291]),
.io_parallelIn_3292(dataIn[3292]),
.io_parallelIn_3293(dataIn[3293]),
.io_parallelIn_3294(dataIn[3294]),
.io_parallelIn_3295(dataIn[3295]),
.io_parallelIn_3296(dataIn[3296]),
.io_parallelIn_3297(dataIn[3297]),
.io_parallelIn_3298(dataIn[3298]),
.io_parallelIn_3299(dataIn[3299]),
.io_parallelIn_3300(dataIn[3300]),
.io_parallelIn_3301(dataIn[3301]),
.io_parallelIn_3302(dataIn[3302]),
.io_parallelIn_3303(dataIn[3303]),
.io_parallelIn_3304(dataIn[3304]),
.io_parallelIn_3305(dataIn[3305]),
.io_parallelIn_3306(dataIn[3306]),
.io_parallelIn_3307(dataIn[3307]),
.io_parallelIn_3308(dataIn[3308]),
.io_parallelIn_3309(dataIn[3309]),
.io_parallelIn_3310(dataIn[3310]),
.io_parallelIn_3311(dataIn[3311]),
.io_parallelIn_3312(dataIn[3312]),
.io_parallelIn_3313(dataIn[3313]),
.io_parallelIn_3314(dataIn[3314]),
.io_parallelIn_3315(dataIn[3315]),
.io_parallelIn_3316(dataIn[3316]),
.io_parallelIn_3317(dataIn[3317]),
.io_parallelIn_3318(dataIn[3318]),
.io_parallelIn_3319(dataIn[3319]),
.io_parallelIn_3320(dataIn[3320]),
.io_parallelIn_3321(dataIn[3321]),
.io_parallelIn_3322(dataIn[3322]),
.io_parallelIn_3323(dataIn[3323]),
.io_parallelIn_3324(dataIn[3324]),
.io_parallelIn_3325(dataIn[3325]),
.io_parallelIn_3326(dataIn[3326]),
.io_parallelIn_3327(dataIn[3327]),
.io_parallelIn_3328(dataIn[3328]),
.io_parallelIn_3329(dataIn[3329]),
.io_parallelIn_3330(dataIn[3330]),
.io_parallelIn_3331(dataIn[3331]),
.io_parallelIn_3332(dataIn[3332]),
.io_parallelIn_3333(dataIn[3333]),
.io_parallelIn_3334(dataIn[3334]),
.io_parallelIn_3335(dataIn[3335]),
.io_parallelIn_3336(dataIn[3336]),
.io_parallelIn_3337(dataIn[3337]),
.io_parallelIn_3338(dataIn[3338]),
.io_parallelIn_3339(dataIn[3339]),
.io_parallelIn_3340(dataIn[3340]),
.io_parallelIn_3341(dataIn[3341]),
.io_parallelIn_3342(dataIn[3342]),
.io_parallelIn_3343(dataIn[3343]),
.io_parallelIn_3344(dataIn[3344]),
.io_parallelIn_3345(dataIn[3345]),
.io_parallelIn_3346(dataIn[3346]),
.io_parallelIn_3347(dataIn[3347]),
.io_parallelIn_3348(dataIn[3348]),
.io_parallelIn_3349(dataIn[3349]),
.io_parallelIn_3350(dataIn[3350]),
.io_parallelIn_3351(dataIn[3351]),
.io_parallelIn_3352(dataIn[3352]),
.io_parallelIn_3353(dataIn[3353]),
.io_parallelIn_3354(dataIn[3354]),
.io_parallelIn_3355(dataIn[3355]),
.io_parallelIn_3356(dataIn[3356]),
.io_parallelIn_3357(dataIn[3357]),
.io_parallelIn_3358(dataIn[3358]),
.io_parallelIn_3359(dataIn[3359]),
.io_parallelIn_3360(dataIn[3360]),
.io_parallelIn_3361(dataIn[3361]),
.io_parallelIn_3362(dataIn[3362]),
.io_parallelIn_3363(dataIn[3363]),
.io_parallelIn_3364(dataIn[3364]),
.io_parallelIn_3365(dataIn[3365]),
.io_parallelIn_3366(dataIn[3366]),
.io_parallelIn_3367(dataIn[3367]),
.io_parallelIn_3368(dataIn[3368]),
.io_parallelIn_3369(dataIn[3369]),
.io_parallelIn_3370(dataIn[3370]),
.io_parallelIn_3371(dataIn[3371]),
.io_parallelIn_3372(dataIn[3372]),
.io_parallelIn_3373(dataIn[3373]),
.io_parallelIn_3374(dataIn[3374]),
.io_parallelIn_3375(dataIn[3375]),
.io_parallelIn_3376(dataIn[3376]),
.io_parallelIn_3377(dataIn[3377]),
.io_parallelIn_3378(dataIn[3378]),
.io_parallelIn_3379(dataIn[3379]),
.io_parallelIn_3380(dataIn[3380]),
.io_parallelIn_3381(dataIn[3381]),
.io_parallelIn_3382(dataIn[3382]),
.io_parallelIn_3383(dataIn[3383]),
.io_parallelIn_3384(dataIn[3384]),
.io_parallelIn_3385(dataIn[3385]),
.io_parallelIn_3386(dataIn[3386]),
.io_parallelIn_3387(dataIn[3387]),
.io_parallelIn_3388(dataIn[3388]),
.io_parallelIn_3389(dataIn[3389]),
.io_parallelIn_3390(dataIn[3390]),
.io_parallelIn_3391(dataIn[3391]),
.io_parallelIn_3392(dataIn[3392]),
.io_parallelIn_3393(dataIn[3393]),
.io_parallelIn_3394(dataIn[3394]),
.io_parallelIn_3395(dataIn[3395]),
.io_parallelIn_3396(dataIn[3396]),
.io_parallelIn_3397(dataIn[3397]),
.io_parallelIn_3398(dataIn[3398]),
.io_parallelIn_3399(dataIn[3399]),
.io_parallelIn_3400(dataIn[3400]),
.io_parallelIn_3401(dataIn[3401]),
.io_parallelIn_3402(dataIn[3402]),
.io_parallelIn_3403(dataIn[3403]),
.io_parallelIn_3404(dataIn[3404]),
.io_parallelIn_3405(dataIn[3405]),
.io_parallelIn_3406(dataIn[3406]),
.io_parallelIn_3407(dataIn[3407]),
.io_parallelIn_3408(dataIn[3408]),
.io_parallelIn_3409(dataIn[3409]),
.io_parallelIn_3410(dataIn[3410]),
.io_parallelIn_3411(dataIn[3411]),
.io_parallelIn_3412(dataIn[3412]),
.io_parallelIn_3413(dataIn[3413]),
.io_parallelIn_3414(dataIn[3414]),
.io_parallelIn_3415(dataIn[3415]),
.io_parallelIn_3416(dataIn[3416]),
.io_parallelIn_3417(dataIn[3417]),
.io_parallelIn_3418(dataIn[3418]),
.io_parallelIn_3419(dataIn[3419]),
.io_parallelIn_3420(dataIn[3420]),
.io_parallelIn_3421(dataIn[3421]),
.io_parallelIn_3422(dataIn[3422]),
.io_parallelIn_3423(dataIn[3423]),
.io_parallelIn_3424(dataIn[3424]),
.io_parallelIn_3425(dataIn[3425]),
.io_parallelIn_3426(dataIn[3426]),
.io_parallelIn_3427(dataIn[3427]),
.io_parallelIn_3428(dataIn[3428]),
.io_parallelIn_3429(dataIn[3429]),
.io_parallelIn_3430(dataIn[3430]),
.io_parallelIn_3431(dataIn[3431]),
.io_parallelIn_3432(dataIn[3432]),
.io_parallelIn_3433(dataIn[3433]),
.io_parallelIn_3434(dataIn[3434]),
.io_parallelIn_3435(dataIn[3435]),
.io_parallelIn_3436(dataIn[3436]),
.io_parallelIn_3437(dataIn[3437]),
.io_parallelIn_3438(dataIn[3438]),
.io_parallelIn_3439(dataIn[3439]),
.io_parallelIn_3440(dataIn[3440]),
.io_parallelIn_3441(dataIn[3441]),
.io_parallelIn_3442(dataIn[3442]),
.io_parallelIn_3443(dataIn[3443]),
.io_parallelIn_3444(dataIn[3444]),
.io_parallelIn_3445(dataIn[3445]),
.io_parallelIn_3446(dataIn[3446]),
.io_parallelIn_3447(dataIn[3447]),
.io_parallelIn_3448(dataIn[3448]),
.io_parallelIn_3449(dataIn[3449]),
.io_parallelIn_3450(dataIn[3450]),
.io_parallelIn_3451(dataIn[3451]),
.io_parallelIn_3452(dataIn[3452]),
.io_parallelIn_3453(dataIn[3453]),
.io_parallelIn_3454(dataIn[3454]),
.io_parallelIn_3455(dataIn[3455]),
.io_parallelIn_3456(dataIn[3456]),
.io_parallelIn_3457(dataIn[3457]),
.io_parallelIn_3458(dataIn[3458]),
.io_parallelIn_3459(dataIn[3459]),
.io_parallelIn_3460(dataIn[3460]),
.io_parallelIn_3461(dataIn[3461]),
.io_parallelIn_3462(dataIn[3462]),
.io_parallelIn_3463(dataIn[3463]),
.io_parallelIn_3464(dataIn[3464]),
.io_parallelIn_3465(dataIn[3465]),
.io_parallelIn_3466(dataIn[3466]),
.io_parallelIn_3467(dataIn[3467]),
.io_parallelIn_3468(dataIn[3468]),
.io_parallelIn_3469(dataIn[3469]),
.io_parallelIn_3470(dataIn[3470]),
.io_parallelIn_3471(dataIn[3471]),
.io_parallelIn_3472(dataIn[3472]),
.io_parallelIn_3473(dataIn[3473]),
.io_parallelIn_3474(dataIn[3474]),
.io_parallelIn_3475(dataIn[3475]),
.io_parallelIn_3476(dataIn[3476]),
.io_parallelIn_3477(dataIn[3477]),
.io_parallelIn_3478(dataIn[3478]),
.io_parallelIn_3479(dataIn[3479]),
.io_parallelIn_3480(dataIn[3480]),
.io_parallelIn_3481(dataIn[3481]),
.io_parallelIn_3482(dataIn[3482]),
.io_parallelIn_3483(dataIn[3483]),
.io_parallelIn_3484(dataIn[3484]),
.io_parallelIn_3485(dataIn[3485]),
.io_parallelIn_3486(dataIn[3486]),
.io_parallelIn_3487(dataIn[3487]),
.io_parallelIn_3488(dataIn[3488]),
.io_parallelIn_3489(dataIn[3489]),
.io_parallelIn_3490(dataIn[3490]),
.io_parallelIn_3491(dataIn[3491]),
.io_parallelIn_3492(dataIn[3492]),
.io_parallelIn_3493(dataIn[3493]),
.io_parallelIn_3494(dataIn[3494]),
.io_parallelIn_3495(dataIn[3495]),
.io_parallelIn_3496(dataIn[3496]),
.io_parallelIn_3497(dataIn[3497]),
.io_parallelIn_3498(dataIn[3498]),
.io_parallelIn_3499(dataIn[3499]),
.io_parallelIn_3500(dataIn[3500]),
.io_parallelIn_3501(dataIn[3501]),
.io_parallelIn_3502(dataIn[3502]),
.io_parallelIn_3503(dataIn[3503]),
.io_parallelIn_3504(dataIn[3504]),
.io_parallelIn_3505(dataIn[3505]),
.io_parallelIn_3506(dataIn[3506]),
.io_parallelIn_3507(dataIn[3507]),
.io_parallelIn_3508(dataIn[3508]),
.io_parallelIn_3509(dataIn[3509]),
.io_parallelIn_3510(dataIn[3510]),
.io_parallelIn_3511(dataIn[3511]),
.io_parallelIn_3512(dataIn[3512]),
.io_parallelIn_3513(dataIn[3513]),
.io_parallelIn_3514(dataIn[3514]),
.io_parallelIn_3515(dataIn[3515]),
.io_parallelIn_3516(dataIn[3516]),
.io_parallelIn_3517(dataIn[3517]),
.io_parallelIn_3518(dataIn[3518]),
.io_parallelIn_3519(dataIn[3519]),
.io_parallelIn_3520(dataIn[3520]),
.io_parallelIn_3521(dataIn[3521]),
.io_parallelIn_3522(dataIn[3522]),
.io_parallelIn_3523(dataIn[3523]),
.io_parallelIn_3524(dataIn[3524]),
.io_parallelIn_3525(dataIn[3525]),
.io_parallelIn_3526(dataIn[3526]),
.io_parallelIn_3527(dataIn[3527]),
.io_parallelIn_3528(dataIn[3528]),
.io_parallelIn_3529(dataIn[3529]),
.io_parallelIn_3530(dataIn[3530]),
.io_parallelIn_3531(dataIn[3531]),
.io_parallelIn_3532(dataIn[3532]),
.io_parallelIn_3533(dataIn[3533]),
.io_parallelIn_3534(dataIn[3534]),
.io_parallelIn_3535(dataIn[3535]),
.io_parallelIn_3536(dataIn[3536]),
.io_parallelIn_3537(dataIn[3537]),
.io_parallelIn_3538(dataIn[3538]),
.io_parallelIn_3539(dataIn[3539]),
.io_parallelIn_3540(dataIn[3540]),
.io_parallelIn_3541(dataIn[3541]),
.io_parallelIn_3542(dataIn[3542]),
.io_parallelIn_3543(dataIn[3543]),
.io_parallelIn_3544(dataIn[3544]),
.io_parallelIn_3545(dataIn[3545]),
.io_parallelIn_3546(dataIn[3546]),
.io_parallelIn_3547(dataIn[3547]),
.io_parallelIn_3548(dataIn[3548]),
.io_parallelIn_3549(dataIn[3549]),
.io_parallelIn_3550(dataIn[3550]),
.io_parallelIn_3551(dataIn[3551]),
.io_parallelIn_3552(dataIn[3552]),
.io_parallelIn_3553(dataIn[3553]),
.io_parallelIn_3554(dataIn[3554]),
.io_parallelIn_3555(dataIn[3555]),
.io_parallelIn_3556(dataIn[3556]),
.io_parallelIn_3557(dataIn[3557]),
.io_parallelIn_3558(dataIn[3558]),
.io_parallelIn_3559(dataIn[3559]),
.io_parallelIn_3560(dataIn[3560]),
.io_parallelIn_3561(dataIn[3561]),
.io_parallelIn_3562(dataIn[3562]),
.io_parallelIn_3563(dataIn[3563]),
.io_parallelIn_3564(dataIn[3564]),
.io_parallelIn_3565(dataIn[3565]),
.io_parallelIn_3566(dataIn[3566]),
.io_parallelIn_3567(dataIn[3567]),
.io_parallelIn_3568(dataIn[3568]),
.io_parallelIn_3569(dataIn[3569]),
.io_parallelIn_3570(dataIn[3570]),
.io_parallelIn_3571(dataIn[3571]),
.io_parallelIn_3572(dataIn[3572]),
.io_parallelIn_3573(dataIn[3573]),
.io_parallelIn_3574(dataIn[3574]),
.io_parallelIn_3575(dataIn[3575]),
.io_parallelIn_3576(dataIn[3576]),
.io_parallelIn_3577(dataIn[3577]),
.io_parallelIn_3578(dataIn[3578]),
.io_parallelIn_3579(dataIn[3579]),
.io_parallelIn_3580(dataIn[3580]),
.io_parallelIn_3581(dataIn[3581]),
.io_parallelIn_3582(dataIn[3582]),
.io_parallelIn_3583(dataIn[3583]),
.io_parallelIn_3584(dataIn[3584]),
.io_parallelIn_3585(dataIn[3585]),
.io_parallelIn_3586(dataIn[3586]),
.io_parallelIn_3587(dataIn[3587]),
.io_parallelIn_3588(dataIn[3588]),
.io_parallelIn_3589(dataIn[3589]),
.io_parallelIn_3590(dataIn[3590]),
.io_parallelIn_3591(dataIn[3591]),
.io_parallelIn_3592(dataIn[3592]),
.io_parallelIn_3593(dataIn[3593]),
.io_parallelIn_3594(dataIn[3594]),
.io_parallelIn_3595(dataIn[3595]),
.io_parallelIn_3596(dataIn[3596]),
.io_parallelIn_3597(dataIn[3597]),
.io_parallelIn_3598(dataIn[3598]),
.io_parallelIn_3599(dataIn[3599]),
.io_parallelIn_3600(dataIn[3600]),
.io_parallelIn_3601(dataIn[3601]),
.io_parallelIn_3602(dataIn[3602]),
.io_parallelIn_3603(dataIn[3603]),
.io_parallelIn_3604(dataIn[3604]),
.io_parallelIn_3605(dataIn[3605]),
.io_parallelIn_3606(dataIn[3606]),
.io_parallelIn_3607(dataIn[3607]),
.io_parallelIn_3608(dataIn[3608]),
.io_parallelIn_3609(dataIn[3609]),
.io_parallelIn_3610(dataIn[3610]),
.io_parallelIn_3611(dataIn[3611]),
.io_parallelIn_3612(dataIn[3612]),
.io_parallelIn_3613(dataIn[3613]),
.io_parallelIn_3614(dataIn[3614]),
.io_parallelIn_3615(dataIn[3615]),
.io_parallelIn_3616(dataIn[3616]),
.io_parallelIn_3617(dataIn[3617]),
.io_parallelIn_3618(dataIn[3618]),
.io_parallelIn_3619(dataIn[3619]),
.io_parallelIn_3620(dataIn[3620]),
.io_parallelIn_3621(dataIn[3621]),
.io_parallelIn_3622(dataIn[3622]),
.io_parallelIn_3623(dataIn[3623]),
.io_parallelIn_3624(dataIn[3624]),
.io_parallelIn_3625(dataIn[3625]),
.io_parallelIn_3626(dataIn[3626]),
.io_parallelIn_3627(dataIn[3627]),
.io_parallelIn_3628(dataIn[3628]),
.io_parallelIn_3629(dataIn[3629]),
.io_parallelIn_3630(dataIn[3630]),
.io_parallelIn_3631(dataIn[3631]),
.io_parallelIn_3632(dataIn[3632]),
.io_parallelIn_3633(dataIn[3633]),
.io_parallelIn_3634(dataIn[3634]),
.io_parallelIn_3635(dataIn[3635]),
.io_parallelIn_3636(dataIn[3636]),
.io_parallelIn_3637(dataIn[3637]),
.io_parallelIn_3638(dataIn[3638]),
.io_parallelIn_3639(dataIn[3639]),
.io_parallelIn_3640(dataIn[3640]),
.io_parallelIn_3641(dataIn[3641]),
.io_parallelIn_3642(dataIn[3642]),
.io_parallelIn_3643(dataIn[3643]),
.io_parallelIn_3644(dataIn[3644]),
.io_parallelIn_3645(dataIn[3645]),
.io_parallelIn_3646(dataIn[3646]),
.io_parallelIn_3647(dataIn[3647]),
.io_parallelIn_3648(dataIn[3648]),
.io_parallelIn_3649(dataIn[3649]),
.io_parallelIn_3650(dataIn[3650]),
.io_parallelIn_3651(dataIn[3651]),
.io_parallelIn_3652(dataIn[3652]),
.io_parallelIn_3653(dataIn[3653]),
.io_parallelIn_3654(dataIn[3654]),
.io_parallelIn_3655(dataIn[3655]),
.io_parallelIn_3656(dataIn[3656]),
.io_parallelIn_3657(dataIn[3657]),
.io_parallelIn_3658(dataIn[3658]),
.io_parallelIn_3659(dataIn[3659]),
.io_parallelIn_3660(dataIn[3660]),
.io_parallelIn_3661(dataIn[3661]),
.io_parallelIn_3662(dataIn[3662]),
.io_parallelIn_3663(dataIn[3663]),
.io_parallelIn_3664(dataIn[3664]),
.io_parallelIn_3665(dataIn[3665]),
.io_parallelIn_3666(dataIn[3666]),
.io_parallelIn_3667(dataIn[3667]),
.io_parallelIn_3668(dataIn[3668]),
.io_parallelIn_3669(dataIn[3669]),
.io_parallelIn_3670(dataIn[3670]),
.io_parallelIn_3671(dataIn[3671]),
.io_parallelIn_3672(dataIn[3672]),
.io_parallelIn_3673(dataIn[3673]),
.io_parallelIn_3674(dataIn[3674]),
.io_parallelIn_3675(dataIn[3675]),
.io_parallelIn_3676(dataIn[3676]),
.io_parallelIn_3677(dataIn[3677]),
.io_parallelIn_3678(dataIn[3678]),
.io_parallelIn_3679(dataIn[3679]),
.io_parallelIn_3680(dataIn[3680]),
.io_parallelIn_3681(dataIn[3681]),
.io_parallelIn_3682(dataIn[3682]),
.io_parallelIn_3683(dataIn[3683]),
.io_parallelIn_3684(dataIn[3684]),
.io_parallelIn_3685(dataIn[3685]),
.io_parallelIn_3686(dataIn[3686]),
.io_parallelIn_3687(dataIn[3687]),
.io_parallelIn_3688(dataIn[3688]),
.io_parallelIn_3689(dataIn[3689]),
.io_parallelIn_3690(dataIn[3690]),
.io_parallelIn_3691(dataIn[3691]),
.io_parallelIn_3692(dataIn[3692]),
.io_parallelIn_3693(dataIn[3693]),
.io_parallelIn_3694(dataIn[3694]),
.io_parallelIn_3695(dataIn[3695]),
.io_parallelIn_3696(dataIn[3696]),
.io_parallelIn_3697(dataIn[3697]),
.io_parallelIn_3698(dataIn[3698]),
.io_parallelIn_3699(dataIn[3699]),
.io_parallelIn_3700(dataIn[3700]),
.io_parallelIn_3701(dataIn[3701]),
.io_parallelIn_3702(dataIn[3702]),
.io_parallelIn_3703(dataIn[3703]),
.io_parallelIn_3704(dataIn[3704]),
.io_parallelIn_3705(dataIn[3705]),
.io_parallelIn_3706(dataIn[3706]),
.io_parallelIn_3707(dataIn[3707]),
.io_parallelIn_3708(dataIn[3708]),
.io_parallelIn_3709(dataIn[3709]),
.io_parallelIn_3710(dataIn[3710]),
.io_parallelIn_3711(dataIn[3711]),
.io_parallelIn_3712(dataIn[3712]),
.io_parallelIn_3713(dataIn[3713]),
.io_parallelIn_3714(dataIn[3714]),
.io_parallelIn_3715(dataIn[3715]),
.io_parallelIn_3716(dataIn[3716]),
.io_parallelIn_3717(dataIn[3717]),
.io_parallelIn_3718(dataIn[3718]),
.io_parallelIn_3719(dataIn[3719]),
.io_parallelIn_3720(dataIn[3720]),
.io_parallelIn_3721(dataIn[3721]),
.io_parallelIn_3722(dataIn[3722]),
.io_parallelIn_3723(dataIn[3723]),
.io_parallelIn_3724(dataIn[3724]),
.io_parallelIn_3725(dataIn[3725]),
.io_parallelIn_3726(dataIn[3726]),
.io_parallelIn_3727(dataIn[3727]),
.io_parallelIn_3728(dataIn[3728]),
.io_parallelIn_3729(dataIn[3729]),
.io_parallelIn_3730(dataIn[3730]),
.io_parallelIn_3731(dataIn[3731]),
.io_parallelIn_3732(dataIn[3732]),
.io_parallelIn_3733(dataIn[3733]),
.io_parallelIn_3734(dataIn[3734]),
.io_parallelIn_3735(dataIn[3735]),
.io_parallelIn_3736(dataIn[3736]),
.io_parallelIn_3737(dataIn[3737]),
.io_parallelIn_3738(dataIn[3738]),
.io_parallelIn_3739(dataIn[3739]),
.io_parallelIn_3740(dataIn[3740]),
.io_parallelIn_3741(dataIn[3741]),
.io_parallelIn_3742(dataIn[3742]),
.io_parallelIn_3743(dataIn[3743]),
.io_parallelIn_3744(dataIn[3744]),
.io_parallelIn_3745(dataIn[3745]),
.io_parallelIn_3746(dataIn[3746]),
.io_parallelIn_3747(dataIn[3747]),
.io_parallelIn_3748(dataIn[3748]),
.io_parallelIn_3749(dataIn[3749]),
.io_parallelIn_3750(dataIn[3750]),
.io_parallelIn_3751(dataIn[3751]),
.io_parallelIn_3752(dataIn[3752]),
.io_parallelIn_3753(dataIn[3753]),
.io_parallelIn_3754(dataIn[3754]),
.io_parallelIn_3755(dataIn[3755]),
.io_parallelIn_3756(dataIn[3756]),
.io_parallelIn_3757(dataIn[3757]),
.io_parallelIn_3758(dataIn[3758]),
.io_parallelIn_3759(dataIn[3759]),
.io_parallelIn_3760(dataIn[3760]),
.io_parallelIn_3761(dataIn[3761]),
.io_parallelIn_3762(dataIn[3762]),
.io_parallelIn_3763(dataIn[3763]),
.io_parallelIn_3764(dataIn[3764]),
.io_parallelIn_3765(dataIn[3765]),
.io_parallelIn_3766(dataIn[3766]),
.io_parallelIn_3767(dataIn[3767]),
.io_parallelIn_3768(dataIn[3768]),
.io_parallelIn_3769(dataIn[3769]),
.io_parallelIn_3770(dataIn[3770]),
.io_parallelIn_3771(dataIn[3771]),
.io_parallelIn_3772(dataIn[3772]),
.io_parallelIn_3773(dataIn[3773]),
.io_parallelIn_3774(dataIn[3774]),
.io_parallelIn_3775(dataIn[3775]),
.io_parallelIn_3776(dataIn[3776]),
.io_parallelIn_3777(dataIn[3777]),
.io_parallelIn_3778(dataIn[3778]),
.io_parallelIn_3779(dataIn[3779]),
.io_parallelIn_3780(dataIn[3780]),
.io_parallelIn_3781(dataIn[3781]),
.io_parallelIn_3782(dataIn[3782]),
.io_parallelIn_3783(dataIn[3783]),
.io_parallelIn_3784(dataIn[3784]),
.io_parallelIn_3785(dataIn[3785]),
.io_parallelIn_3786(dataIn[3786]),
.io_parallelIn_3787(dataIn[3787]),
.io_parallelIn_3788(dataIn[3788]),
.io_parallelIn_3789(dataIn[3789]),
.io_parallelIn_3790(dataIn[3790]),
.io_parallelIn_3791(dataIn[3791]),
.io_parallelIn_3792(dataIn[3792]),
.io_parallelIn_3793(dataIn[3793]),
.io_parallelIn_3794(dataIn[3794]),
.io_parallelIn_3795(dataIn[3795]),
.io_parallelIn_3796(dataIn[3796]),
.io_parallelIn_3797(dataIn[3797]),
.io_parallelIn_3798(dataIn[3798]),
.io_parallelIn_3799(dataIn[3799]),
.io_parallelIn_3800(dataIn[3800]),
.io_parallelIn_3801(dataIn[3801]),
.io_parallelIn_3802(dataIn[3802]),
.io_parallelIn_3803(dataIn[3803]),
.io_parallelIn_3804(dataIn[3804]),
.io_parallelIn_3805(dataIn[3805]),
.io_parallelIn_3806(dataIn[3806]),
.io_parallelIn_3807(dataIn[3807]),
.io_parallelIn_3808(dataIn[3808]),
.io_parallelIn_3809(dataIn[3809]),
.io_parallelIn_3810(dataIn[3810]),
.io_parallelIn_3811(dataIn[3811]),
.io_parallelIn_3812(dataIn[3812]),
.io_parallelIn_3813(dataIn[3813]),
.io_parallelIn_3814(dataIn[3814]),
.io_parallelIn_3815(dataIn[3815]),
.io_parallelIn_3816(dataIn[3816]),
.io_parallelIn_3817(dataIn[3817]),
.io_parallelIn_3818(dataIn[3818]),
.io_parallelIn_3819(dataIn[3819]),
.io_parallelIn_3820(dataIn[3820]),
.io_parallelIn_3821(dataIn[3821]),
.io_parallelIn_3822(dataIn[3822]),
.io_parallelIn_3823(dataIn[3823]),
.io_parallelIn_3824(dataIn[3824]),
.io_parallelIn_3825(dataIn[3825]),
.io_parallelIn_3826(dataIn[3826]),
.io_parallelIn_3827(dataIn[3827]),
.io_parallelIn_3828(dataIn[3828]),
.io_parallelIn_3829(dataIn[3829]),
.io_parallelIn_3830(dataIn[3830]),
.io_parallelIn_3831(dataIn[3831]),
.io_parallelIn_3832(dataIn[3832]),
.io_parallelIn_3833(dataIn[3833]),
.io_parallelIn_3834(dataIn[3834]),
.io_parallelIn_3835(dataIn[3835]),
.io_parallelIn_3836(dataIn[3836]),
.io_parallelIn_3837(dataIn[3837]),
.io_parallelIn_3838(dataIn[3838]),
.io_parallelIn_3839(dataIn[3839]),
.io_parallelIn_3840(dataIn[3840]),
.io_parallelIn_3841(dataIn[3841]),
.io_parallelIn_3842(dataIn[3842]),
.io_parallelIn_3843(dataIn[3843]),
.io_parallelIn_3844(dataIn[3844]),
.io_parallelIn_3845(dataIn[3845]),
.io_parallelIn_3846(dataIn[3846]),
.io_parallelIn_3847(dataIn[3847]),
.io_parallelIn_3848(dataIn[3848]),
.io_parallelIn_3849(dataIn[3849]),
.io_parallelIn_3850(dataIn[3850]),
.io_parallelIn_3851(dataIn[3851]),
.io_parallelIn_3852(dataIn[3852]),
.io_parallelIn_3853(dataIn[3853]),
.io_parallelIn_3854(dataIn[3854]),
.io_parallelIn_3855(dataIn[3855]),
.io_parallelIn_3856(dataIn[3856]),
.io_parallelIn_3857(dataIn[3857]),
.io_parallelIn_3858(dataIn[3858]),
.io_parallelIn_3859(dataIn[3859]),
.io_parallelIn_3860(dataIn[3860]),
.io_parallelIn_3861(dataIn[3861]),
.io_parallelIn_3862(dataIn[3862]),
.io_parallelIn_3863(dataIn[3863]),
.io_parallelIn_3864(dataIn[3864]),
.io_parallelIn_3865(dataIn[3865]),
.io_parallelIn_3866(dataIn[3866]),
.io_parallelIn_3867(dataIn[3867]),
.io_parallelIn_3868(dataIn[3868]),
.io_parallelIn_3869(dataIn[3869]),
.io_parallelIn_3870(dataIn[3870]),
.io_parallelIn_3871(dataIn[3871]),
.io_parallelIn_3872(dataIn[3872]),
.io_parallelIn_3873(dataIn[3873]),
.io_parallelIn_3874(dataIn[3874]),
.io_parallelIn_3875(dataIn[3875]),
.io_parallelIn_3876(dataIn[3876]),
.io_parallelIn_3877(dataIn[3877]),
.io_parallelIn_3878(dataIn[3878]),
.io_parallelIn_3879(dataIn[3879]),
.io_parallelIn_3880(dataIn[3880]),
.io_parallelIn_3881(dataIn[3881]),
.io_parallelIn_3882(dataIn[3882]),
.io_parallelIn_3883(dataIn[3883]),
.io_parallelIn_3884(dataIn[3884]),
.io_parallelIn_3885(dataIn[3885]),
.io_parallelIn_3886(dataIn[3886]),
.io_parallelIn_3887(dataIn[3887]),
.io_parallelIn_3888(dataIn[3888]),
.io_parallelIn_3889(dataIn[3889]),
.io_parallelIn_3890(dataIn[3890]),
.io_parallelIn_3891(dataIn[3891]),
.io_parallelIn_3892(dataIn[3892]),
.io_parallelIn_3893(dataIn[3893]),
.io_parallelIn_3894(dataIn[3894]),
.io_parallelIn_3895(dataIn[3895]),
.io_parallelIn_3896(dataIn[3896]),
.io_parallelIn_3897(dataIn[3897]),
.io_parallelIn_3898(dataIn[3898]),
.io_parallelIn_3899(dataIn[3899]),
.io_parallelIn_3900(dataIn[3900]),
.io_parallelIn_3901(dataIn[3901]),
.io_parallelIn_3902(dataIn[3902]),
.io_parallelIn_3903(dataIn[3903]),
.io_parallelIn_3904(dataIn[3904]),
.io_parallelIn_3905(dataIn[3905]),
.io_parallelIn_3906(dataIn[3906]),
.io_parallelIn_3907(dataIn[3907]),
.io_parallelIn_3908(dataIn[3908]),
.io_parallelIn_3909(dataIn[3909]),
.io_parallelIn_3910(dataIn[3910]),
.io_parallelIn_3911(dataIn[3911]),
.io_parallelIn_3912(dataIn[3912]),
.io_parallelIn_3913(dataIn[3913]),
.io_parallelIn_3914(dataIn[3914]),
.io_parallelIn_3915(dataIn[3915]),
.io_parallelIn_3916(dataIn[3916]),
.io_parallelIn_3917(dataIn[3917]),
.io_parallelIn_3918(dataIn[3918]),
.io_parallelIn_3919(dataIn[3919]),
.io_parallelIn_3920(dataIn[3920]),
.io_parallelIn_3921(dataIn[3921]),
.io_parallelIn_3922(dataIn[3922]),
.io_parallelIn_3923(dataIn[3923]),
.io_parallelIn_3924(dataIn[3924]),
.io_parallelIn_3925(dataIn[3925]),
.io_parallelIn_3926(dataIn[3926]),
.io_parallelIn_3927(dataIn[3927]),
.io_parallelIn_3928(dataIn[3928]),
.io_parallelIn_3929(dataIn[3929]),
.io_parallelIn_3930(dataIn[3930]),
.io_parallelIn_3931(dataIn[3931]),
.io_parallelIn_3932(dataIn[3932]),
.io_parallelIn_3933(dataIn[3933]),
.io_parallelIn_3934(dataIn[3934]),
.io_parallelIn_3935(dataIn[3935]),
.io_parallelIn_3936(dataIn[3936]),
.io_parallelIn_3937(dataIn[3937]),
.io_parallelIn_3938(dataIn[3938]),
.io_parallelIn_3939(dataIn[3939]),
.io_parallelIn_3940(dataIn[3940]),
.io_parallelIn_3941(dataIn[3941]),
.io_parallelIn_3942(dataIn[3942]),
.io_parallelIn_3943(dataIn[3943]),
.io_parallelIn_3944(dataIn[3944]),
.io_parallelIn_3945(dataIn[3945]),
.io_parallelIn_3946(dataIn[3946]),
.io_parallelIn_3947(dataIn[3947]),
.io_parallelIn_3948(dataIn[3948]),
.io_parallelIn_3949(dataIn[3949]),
.io_parallelIn_3950(dataIn[3950]),
.io_parallelIn_3951(dataIn[3951]),
.io_parallelIn_3952(dataIn[3952]),
.io_parallelIn_3953(dataIn[3953]),
.io_parallelIn_3954(dataIn[3954]),
.io_parallelIn_3955(dataIn[3955]),
.io_parallelIn_3956(dataIn[3956]),
.io_parallelIn_3957(dataIn[3957]),
.io_parallelIn_3958(dataIn[3958]),
.io_parallelIn_3959(dataIn[3959]),
.io_parallelIn_3960(dataIn[3960]),
.io_parallelIn_3961(dataIn[3961]),
.io_parallelIn_3962(dataIn[3962]),
.io_parallelIn_3963(dataIn[3963]),
.io_parallelIn_3964(dataIn[3964]),
.io_parallelIn_3965(dataIn[3965]),
.io_parallelIn_3966(dataIn[3966]),
.io_parallelIn_3967(dataIn[3967]),
.io_parallelIn_3968(dataIn[3968]),
.io_parallelIn_3969(dataIn[3969]),
.io_parallelIn_3970(dataIn[3970]),
.io_parallelIn_3971(dataIn[3971]),
.io_parallelIn_3972(dataIn[3972]),
.io_parallelIn_3973(dataIn[3973]),
.io_parallelIn_3974(dataIn[3974]),
.io_parallelIn_3975(dataIn[3975]),
.io_parallelIn_3976(dataIn[3976]),
.io_parallelIn_3977(dataIn[3977]),
.io_parallelIn_3978(dataIn[3978]),
.io_parallelIn_3979(dataIn[3979]),
.io_parallelIn_3980(dataIn[3980]),
.io_parallelIn_3981(dataIn[3981]),
.io_parallelIn_3982(dataIn[3982]),
.io_parallelIn_3983(dataIn[3983]),
.io_parallelIn_3984(dataIn[3984]),
.io_parallelIn_3985(dataIn[3985]),
.io_parallelIn_3986(dataIn[3986]),
.io_parallelIn_3987(dataIn[3987]),
.io_parallelIn_3988(dataIn[3988]),
.io_parallelIn_3989(dataIn[3989]),
.io_parallelIn_3990(dataIn[3990]),
.io_parallelIn_3991(dataIn[3991]),
.io_parallelIn_3992(dataIn[3992]),
.io_parallelIn_3993(dataIn[3993]),
.io_parallelIn_3994(dataIn[3994]),
.io_parallelIn_3995(dataIn[3995]),
.io_parallelIn_3996(dataIn[3996]),
.io_parallelIn_3997(dataIn[3997]),
.io_parallelIn_3998(dataIn[3998]),
.io_parallelIn_3999(dataIn[3999]),
.io_parallelIn_4000(dataIn[4000]),
.io_parallelIn_4001(dataIn[4001]),
.io_parallelIn_4002(dataIn[4002]),
.io_parallelIn_4003(dataIn[4003]),
.io_parallelIn_4004(dataIn[4004]),
.io_parallelIn_4005(dataIn[4005]),
.io_parallelIn_4006(dataIn[4006]),
.io_parallelIn_4007(dataIn[4007]),
.io_parallelIn_4008(dataIn[4008]),
.io_parallelIn_4009(dataIn[4009]),
.io_parallelIn_4010(dataIn[4010]),
.io_parallelIn_4011(dataIn[4011]),
.io_parallelIn_4012(dataIn[4012]),
.io_parallelIn_4013(dataIn[4013]),
.io_parallelIn_4014(dataIn[4014]),
.io_parallelIn_4015(dataIn[4015]),
.io_parallelIn_4016(dataIn[4016]),
.io_parallelIn_4017(dataIn[4017]),
.io_parallelIn_4018(dataIn[4018]),
.io_parallelIn_4019(dataIn[4019]),
.io_parallelIn_4020(dataIn[4020]),
.io_parallelIn_4021(dataIn[4021]),
.io_parallelIn_4022(dataIn[4022]),
.io_parallelIn_4023(dataIn[4023]),
.io_parallelIn_4024(dataIn[4024]),
.io_parallelIn_4025(dataIn[4025]),
.io_parallelIn_4026(dataIn[4026]),
.io_parallelIn_4027(dataIn[4027]),
.io_parallelIn_4028(dataIn[4028]),
.io_parallelIn_4029(dataIn[4029]),
.io_parallelIn_4030(dataIn[4030]),
.io_parallelIn_4031(dataIn[4031]),
.io_parallelIn_4032(dataIn[4032]),
.io_parallelIn_4033(dataIn[4033]),
.io_parallelIn_4034(dataIn[4034]),
.io_parallelIn_4035(dataIn[4035]),
.io_parallelIn_4036(dataIn[4036]),
.io_parallelIn_4037(dataIn[4037]),
.io_parallelIn_4038(dataIn[4038]),
.io_parallelIn_4039(dataIn[4039]),
.io_parallelIn_4040(dataIn[4040]),
.io_parallelIn_4041(dataIn[4041]),
.io_parallelIn_4042(dataIn[4042]),
.io_parallelIn_4043(dataIn[4043]),
.io_parallelIn_4044(dataIn[4044]),
.io_parallelIn_4045(dataIn[4045]),
.io_parallelIn_4046(dataIn[4046]),
.io_parallelIn_4047(dataIn[4047]),
.io_parallelIn_4048(dataIn[4048]),
.io_parallelIn_4049(dataIn[4049]),
.io_parallelIn_4050(dataIn[4050]),
.io_parallelIn_4051(dataIn[4051]),
.io_parallelIn_4052(dataIn[4052]),
.io_parallelIn_4053(dataIn[4053]),
.io_parallelIn_4054(dataIn[4054]),
.io_parallelIn_4055(dataIn[4055]),
.io_parallelIn_4056(dataIn[4056]),
.io_parallelIn_4057(dataIn[4057]),
.io_parallelIn_4058(dataIn[4058]),
.io_parallelIn_4059(dataIn[4059]),
.io_parallelIn_4060(dataIn[4060]),
.io_parallelIn_4061(dataIn[4061]),
.io_parallelIn_4062(dataIn[4062]),
.io_parallelIn_4063(dataIn[4063]),
.io_parallelIn_4064(dataIn[4064]),
.io_parallelIn_4065(dataIn[4065]),
.io_parallelIn_4066(dataIn[4066]),
.io_parallelIn_4067(dataIn[4067]),
.io_parallelIn_4068(dataIn[4068]),
.io_parallelIn_4069(dataIn[4069]),
.io_parallelIn_4070(dataIn[4070]),
.io_parallelIn_4071(dataIn[4071]),
.io_parallelIn_4072(dataIn[4072]),
.io_parallelIn_4073(dataIn[4073]),
.io_parallelIn_4074(dataIn[4074]),
.io_parallelIn_4075(dataIn[4075]),
.io_parallelIn_4076(dataIn[4076]),
.io_parallelIn_4077(dataIn[4077]),
.io_parallelIn_4078(dataIn[4078]),
.io_parallelIn_4079(dataIn[4079]),
.io_parallelIn_4080(dataIn[4080]),
.io_parallelIn_4081(dataIn[4081]),
.io_parallelIn_4082(dataIn[4082]),
.io_parallelIn_4083(dataIn[4083]),
.io_parallelIn_4084(dataIn[4084]),
.io_parallelIn_4085(dataIn[4085]),
.io_parallelIn_4086(dataIn[4086]),
.io_parallelIn_4087(dataIn[4087]),
.io_parallelIn_4088(dataIn[4088]),
.io_parallelIn_4089(dataIn[4089]),
.io_parallelIn_4090(dataIn[4090]),
.io_parallelIn_4091(dataIn[4091]),
.io_parallelIn_4092(dataIn[4092]),
.io_parallelIn_4093(dataIn[4093]),
.io_parallelIn_4094(dataIn[4094]),
.io_parallelIn_4095(dataIn[4095]),
.io_parallelOut_0(dataOut[0]),
.io_parallelOut_1(dataOut[1]),
.io_parallelOut_2(dataOut[2]),
.io_parallelOut_3(dataOut[3]),
.io_parallelOut_4(dataOut[4]),
.io_parallelOut_5(dataOut[5]),
.io_parallelOut_6(dataOut[6]),
.io_parallelOut_7(dataOut[7]),
.io_parallelOut_8(dataOut[8]),
.io_parallelOut_9(dataOut[9]),
.io_parallelOut_10(dataOut[10]),
.io_parallelOut_11(dataOut[11]),
.io_parallelOut_12(dataOut[12]),
.io_parallelOut_13(dataOut[13]),
.io_parallelOut_14(dataOut[14]),
.io_parallelOut_15(dataOut[15]),
.io_parallelOut_16(dataOut[16]),
.io_parallelOut_17(dataOut[17]),
.io_parallelOut_18(dataOut[18]),
.io_parallelOut_19(dataOut[19]),
.io_parallelOut_20(dataOut[20]),
.io_parallelOut_21(dataOut[21]),
.io_parallelOut_22(dataOut[22]),
.io_parallelOut_23(dataOut[23]),
.io_parallelOut_24(dataOut[24]),
.io_parallelOut_25(dataOut[25]),
.io_parallelOut_26(dataOut[26]),
.io_parallelOut_27(dataOut[27]),
.io_parallelOut_28(dataOut[28]),
.io_parallelOut_29(dataOut[29]),
.io_parallelOut_30(dataOut[30]),
.io_parallelOut_31(dataOut[31]),
.io_parallelOut_32(dataOut[32]),
.io_parallelOut_33(dataOut[33]),
.io_parallelOut_34(dataOut[34]),
.io_parallelOut_35(dataOut[35]),
.io_parallelOut_36(dataOut[36]),
.io_parallelOut_37(dataOut[37]),
.io_parallelOut_38(dataOut[38]),
.io_parallelOut_39(dataOut[39]),
.io_parallelOut_40(dataOut[40]),
.io_parallelOut_41(dataOut[41]),
.io_parallelOut_42(dataOut[42]),
.io_parallelOut_43(dataOut[43]),
.io_parallelOut_44(dataOut[44]),
.io_parallelOut_45(dataOut[45]),
.io_parallelOut_46(dataOut[46]),
.io_parallelOut_47(dataOut[47]),
.io_parallelOut_48(dataOut[48]),
.io_parallelOut_49(dataOut[49]),
.io_parallelOut_50(dataOut[50]),
.io_parallelOut_51(dataOut[51]),
.io_parallelOut_52(dataOut[52]),
.io_parallelOut_53(dataOut[53]),
.io_parallelOut_54(dataOut[54]),
.io_parallelOut_55(dataOut[55]),
.io_parallelOut_56(dataOut[56]),
.io_parallelOut_57(dataOut[57]),
.io_parallelOut_58(dataOut[58]),
.io_parallelOut_59(dataOut[59]),
.io_parallelOut_60(dataOut[60]),
.io_parallelOut_61(dataOut[61]),
.io_parallelOut_62(dataOut[62]),
.io_parallelOut_63(dataOut[63]),
.io_parallelOut_64(dataOut[64]),
.io_parallelOut_65(dataOut[65]),
.io_parallelOut_66(dataOut[66]),
.io_parallelOut_67(dataOut[67]),
.io_parallelOut_68(dataOut[68]),
.io_parallelOut_69(dataOut[69]),
.io_parallelOut_70(dataOut[70]),
.io_parallelOut_71(dataOut[71]),
.io_parallelOut_72(dataOut[72]),
.io_parallelOut_73(dataOut[73]),
.io_parallelOut_74(dataOut[74]),
.io_parallelOut_75(dataOut[75]),
.io_parallelOut_76(dataOut[76]),
.io_parallelOut_77(dataOut[77]),
.io_parallelOut_78(dataOut[78]),
.io_parallelOut_79(dataOut[79]),
.io_parallelOut_80(dataOut[80]),
.io_parallelOut_81(dataOut[81]),
.io_parallelOut_82(dataOut[82]),
.io_parallelOut_83(dataOut[83]),
.io_parallelOut_84(dataOut[84]),
.io_parallelOut_85(dataOut[85]),
.io_parallelOut_86(dataOut[86]),
.io_parallelOut_87(dataOut[87]),
.io_parallelOut_88(dataOut[88]),
.io_parallelOut_89(dataOut[89]),
.io_parallelOut_90(dataOut[90]),
.io_parallelOut_91(dataOut[91]),
.io_parallelOut_92(dataOut[92]),
.io_parallelOut_93(dataOut[93]),
.io_parallelOut_94(dataOut[94]),
.io_parallelOut_95(dataOut[95]),
.io_parallelOut_96(dataOut[96]),
.io_parallelOut_97(dataOut[97]),
.io_parallelOut_98(dataOut[98]),
.io_parallelOut_99(dataOut[99]),
.io_parallelOut_100(dataOut[100]),
.io_parallelOut_101(dataOut[101]),
.io_parallelOut_102(dataOut[102]),
.io_parallelOut_103(dataOut[103]),
.io_parallelOut_104(dataOut[104]),
.io_parallelOut_105(dataOut[105]),
.io_parallelOut_106(dataOut[106]),
.io_parallelOut_107(dataOut[107]),
.io_parallelOut_108(dataOut[108]),
.io_parallelOut_109(dataOut[109]),
.io_parallelOut_110(dataOut[110]),
.io_parallelOut_111(dataOut[111]),
.io_parallelOut_112(dataOut[112]),
.io_parallelOut_113(dataOut[113]),
.io_parallelOut_114(dataOut[114]),
.io_parallelOut_115(dataOut[115]),
.io_parallelOut_116(dataOut[116]),
.io_parallelOut_117(dataOut[117]),
.io_parallelOut_118(dataOut[118]),
.io_parallelOut_119(dataOut[119]),
.io_parallelOut_120(dataOut[120]),
.io_parallelOut_121(dataOut[121]),
.io_parallelOut_122(dataOut[122]),
.io_parallelOut_123(dataOut[123]),
.io_parallelOut_124(dataOut[124]),
.io_parallelOut_125(dataOut[125]),
.io_parallelOut_126(dataOut[126]),
.io_parallelOut_127(dataOut[127]),
.io_parallelOut_128(dataOut[128]),
.io_parallelOut_129(dataOut[129]),
.io_parallelOut_130(dataOut[130]),
.io_parallelOut_131(dataOut[131]),
.io_parallelOut_132(dataOut[132]),
.io_parallelOut_133(dataOut[133]),
.io_parallelOut_134(dataOut[134]),
.io_parallelOut_135(dataOut[135]),
.io_parallelOut_136(dataOut[136]),
.io_parallelOut_137(dataOut[137]),
.io_parallelOut_138(dataOut[138]),
.io_parallelOut_139(dataOut[139]),
.io_parallelOut_140(dataOut[140]),
.io_parallelOut_141(dataOut[141]),
.io_parallelOut_142(dataOut[142]),
.io_parallelOut_143(dataOut[143]),
.io_parallelOut_144(dataOut[144]),
.io_parallelOut_145(dataOut[145]),
.io_parallelOut_146(dataOut[146]),
.io_parallelOut_147(dataOut[147]),
.io_parallelOut_148(dataOut[148]),
.io_parallelOut_149(dataOut[149]),
.io_parallelOut_150(dataOut[150]),
.io_parallelOut_151(dataOut[151]),
.io_parallelOut_152(dataOut[152]),
.io_parallelOut_153(dataOut[153]),
.io_parallelOut_154(dataOut[154]),
.io_parallelOut_155(dataOut[155]),
.io_parallelOut_156(dataOut[156]),
.io_parallelOut_157(dataOut[157]),
.io_parallelOut_158(dataOut[158]),
.io_parallelOut_159(dataOut[159]),
.io_parallelOut_160(dataOut[160]),
.io_parallelOut_161(dataOut[161]),
.io_parallelOut_162(dataOut[162]),
.io_parallelOut_163(dataOut[163]),
.io_parallelOut_164(dataOut[164]),
.io_parallelOut_165(dataOut[165]),
.io_parallelOut_166(dataOut[166]),
.io_parallelOut_167(dataOut[167]),
.io_parallelOut_168(dataOut[168]),
.io_parallelOut_169(dataOut[169]),
.io_parallelOut_170(dataOut[170]),
.io_parallelOut_171(dataOut[171]),
.io_parallelOut_172(dataOut[172]),
.io_parallelOut_173(dataOut[173]),
.io_parallelOut_174(dataOut[174]),
.io_parallelOut_175(dataOut[175]),
.io_parallelOut_176(dataOut[176]),
.io_parallelOut_177(dataOut[177]),
.io_parallelOut_178(dataOut[178]),
.io_parallelOut_179(dataOut[179]),
.io_parallelOut_180(dataOut[180]),
.io_parallelOut_181(dataOut[181]),
.io_parallelOut_182(dataOut[182]),
.io_parallelOut_183(dataOut[183]),
.io_parallelOut_184(dataOut[184]),
.io_parallelOut_185(dataOut[185]),
.io_parallelOut_186(dataOut[186]),
.io_parallelOut_187(dataOut[187]),
.io_parallelOut_188(dataOut[188]),
.io_parallelOut_189(dataOut[189]),
.io_parallelOut_190(dataOut[190]),
.io_parallelOut_191(dataOut[191]),
.io_parallelOut_192(dataOut[192]),
.io_parallelOut_193(dataOut[193]),
.io_parallelOut_194(dataOut[194]),
.io_parallelOut_195(dataOut[195]),
.io_parallelOut_196(dataOut[196]),
.io_parallelOut_197(dataOut[197]),
.io_parallelOut_198(dataOut[198]),
.io_parallelOut_199(dataOut[199]),
.io_parallelOut_200(dataOut[200]),
.io_parallelOut_201(dataOut[201]),
.io_parallelOut_202(dataOut[202]),
.io_parallelOut_203(dataOut[203]),
.io_parallelOut_204(dataOut[204]),
.io_parallelOut_205(dataOut[205]),
.io_parallelOut_206(dataOut[206]),
.io_parallelOut_207(dataOut[207]),
.io_parallelOut_208(dataOut[208]),
.io_parallelOut_209(dataOut[209]),
.io_parallelOut_210(dataOut[210]),
.io_parallelOut_211(dataOut[211]),
.io_parallelOut_212(dataOut[212]),
.io_parallelOut_213(dataOut[213]),
.io_parallelOut_214(dataOut[214]),
.io_parallelOut_215(dataOut[215]),
.io_parallelOut_216(dataOut[216]),
.io_parallelOut_217(dataOut[217]),
.io_parallelOut_218(dataOut[218]),
.io_parallelOut_219(dataOut[219]),
.io_parallelOut_220(dataOut[220]),
.io_parallelOut_221(dataOut[221]),
.io_parallelOut_222(dataOut[222]),
.io_parallelOut_223(dataOut[223]),
.io_parallelOut_224(dataOut[224]),
.io_parallelOut_225(dataOut[225]),
.io_parallelOut_226(dataOut[226]),
.io_parallelOut_227(dataOut[227]),
.io_parallelOut_228(dataOut[228]),
.io_parallelOut_229(dataOut[229]),
.io_parallelOut_230(dataOut[230]),
.io_parallelOut_231(dataOut[231]),
.io_parallelOut_232(dataOut[232]),
.io_parallelOut_233(dataOut[233]),
.io_parallelOut_234(dataOut[234]),
.io_parallelOut_235(dataOut[235]),
.io_parallelOut_236(dataOut[236]),
.io_parallelOut_237(dataOut[237]),
.io_parallelOut_238(dataOut[238]),
.io_parallelOut_239(dataOut[239]),
.io_parallelOut_240(dataOut[240]),
.io_parallelOut_241(dataOut[241]),
.io_parallelOut_242(dataOut[242]),
.io_parallelOut_243(dataOut[243]),
.io_parallelOut_244(dataOut[244]),
.io_parallelOut_245(dataOut[245]),
.io_parallelOut_246(dataOut[246]),
.io_parallelOut_247(dataOut[247]),
.io_parallelOut_248(dataOut[248]),
.io_parallelOut_249(dataOut[249]),
.io_parallelOut_250(dataOut[250]),
.io_parallelOut_251(dataOut[251]),
.io_parallelOut_252(dataOut[252]),
.io_parallelOut_253(dataOut[253]),
.io_parallelOut_254(dataOut[254]),
.io_parallelOut_255(dataOut[255]),
.io_parallelOut_256(dataOut[256]),
.io_parallelOut_257(dataOut[257]),
.io_parallelOut_258(dataOut[258]),
.io_parallelOut_259(dataOut[259]),
.io_parallelOut_260(dataOut[260]),
.io_parallelOut_261(dataOut[261]),
.io_parallelOut_262(dataOut[262]),
.io_parallelOut_263(dataOut[263]),
.io_parallelOut_264(dataOut[264]),
.io_parallelOut_265(dataOut[265]),
.io_parallelOut_266(dataOut[266]),
.io_parallelOut_267(dataOut[267]),
.io_parallelOut_268(dataOut[268]),
.io_parallelOut_269(dataOut[269]),
.io_parallelOut_270(dataOut[270]),
.io_parallelOut_271(dataOut[271]),
.io_parallelOut_272(dataOut[272]),
.io_parallelOut_273(dataOut[273]),
.io_parallelOut_274(dataOut[274]),
.io_parallelOut_275(dataOut[275]),
.io_parallelOut_276(dataOut[276]),
.io_parallelOut_277(dataOut[277]),
.io_parallelOut_278(dataOut[278]),
.io_parallelOut_279(dataOut[279]),
.io_parallelOut_280(dataOut[280]),
.io_parallelOut_281(dataOut[281]),
.io_parallelOut_282(dataOut[282]),
.io_parallelOut_283(dataOut[283]),
.io_parallelOut_284(dataOut[284]),
.io_parallelOut_285(dataOut[285]),
.io_parallelOut_286(dataOut[286]),
.io_parallelOut_287(dataOut[287]),
.io_parallelOut_288(dataOut[288]),
.io_parallelOut_289(dataOut[289]),
.io_parallelOut_290(dataOut[290]),
.io_parallelOut_291(dataOut[291]),
.io_parallelOut_292(dataOut[292]),
.io_parallelOut_293(dataOut[293]),
.io_parallelOut_294(dataOut[294]),
.io_parallelOut_295(dataOut[295]),
.io_parallelOut_296(dataOut[296]),
.io_parallelOut_297(dataOut[297]),
.io_parallelOut_298(dataOut[298]),
.io_parallelOut_299(dataOut[299]),
.io_parallelOut_300(dataOut[300]),
.io_parallelOut_301(dataOut[301]),
.io_parallelOut_302(dataOut[302]),
.io_parallelOut_303(dataOut[303]),
.io_parallelOut_304(dataOut[304]),
.io_parallelOut_305(dataOut[305]),
.io_parallelOut_306(dataOut[306]),
.io_parallelOut_307(dataOut[307]),
.io_parallelOut_308(dataOut[308]),
.io_parallelOut_309(dataOut[309]),
.io_parallelOut_310(dataOut[310]),
.io_parallelOut_311(dataOut[311]),
.io_parallelOut_312(dataOut[312]),
.io_parallelOut_313(dataOut[313]),
.io_parallelOut_314(dataOut[314]),
.io_parallelOut_315(dataOut[315]),
.io_parallelOut_316(dataOut[316]),
.io_parallelOut_317(dataOut[317]),
.io_parallelOut_318(dataOut[318]),
.io_parallelOut_319(dataOut[319]),
.io_parallelOut_320(dataOut[320]),
.io_parallelOut_321(dataOut[321]),
.io_parallelOut_322(dataOut[322]),
.io_parallelOut_323(dataOut[323]),
.io_parallelOut_324(dataOut[324]),
.io_parallelOut_325(dataOut[325]),
.io_parallelOut_326(dataOut[326]),
.io_parallelOut_327(dataOut[327]),
.io_parallelOut_328(dataOut[328]),
.io_parallelOut_329(dataOut[329]),
.io_parallelOut_330(dataOut[330]),
.io_parallelOut_331(dataOut[331]),
.io_parallelOut_332(dataOut[332]),
.io_parallelOut_333(dataOut[333]),
.io_parallelOut_334(dataOut[334]),
.io_parallelOut_335(dataOut[335]),
.io_parallelOut_336(dataOut[336]),
.io_parallelOut_337(dataOut[337]),
.io_parallelOut_338(dataOut[338]),
.io_parallelOut_339(dataOut[339]),
.io_parallelOut_340(dataOut[340]),
.io_parallelOut_341(dataOut[341]),
.io_parallelOut_342(dataOut[342]),
.io_parallelOut_343(dataOut[343]),
.io_parallelOut_344(dataOut[344]),
.io_parallelOut_345(dataOut[345]),
.io_parallelOut_346(dataOut[346]),
.io_parallelOut_347(dataOut[347]),
.io_parallelOut_348(dataOut[348]),
.io_parallelOut_349(dataOut[349]),
.io_parallelOut_350(dataOut[350]),
.io_parallelOut_351(dataOut[351]),
.io_parallelOut_352(dataOut[352]),
.io_parallelOut_353(dataOut[353]),
.io_parallelOut_354(dataOut[354]),
.io_parallelOut_355(dataOut[355]),
.io_parallelOut_356(dataOut[356]),
.io_parallelOut_357(dataOut[357]),
.io_parallelOut_358(dataOut[358]),
.io_parallelOut_359(dataOut[359]),
.io_parallelOut_360(dataOut[360]),
.io_parallelOut_361(dataOut[361]),
.io_parallelOut_362(dataOut[362]),
.io_parallelOut_363(dataOut[363]),
.io_parallelOut_364(dataOut[364]),
.io_parallelOut_365(dataOut[365]),
.io_parallelOut_366(dataOut[366]),
.io_parallelOut_367(dataOut[367]),
.io_parallelOut_368(dataOut[368]),
.io_parallelOut_369(dataOut[369]),
.io_parallelOut_370(dataOut[370]),
.io_parallelOut_371(dataOut[371]),
.io_parallelOut_372(dataOut[372]),
.io_parallelOut_373(dataOut[373]),
.io_parallelOut_374(dataOut[374]),
.io_parallelOut_375(dataOut[375]),
.io_parallelOut_376(dataOut[376]),
.io_parallelOut_377(dataOut[377]),
.io_parallelOut_378(dataOut[378]),
.io_parallelOut_379(dataOut[379]),
.io_parallelOut_380(dataOut[380]),
.io_parallelOut_381(dataOut[381]),
.io_parallelOut_382(dataOut[382]),
.io_parallelOut_383(dataOut[383]),
.io_parallelOut_384(dataOut[384]),
.io_parallelOut_385(dataOut[385]),
.io_parallelOut_386(dataOut[386]),
.io_parallelOut_387(dataOut[387]),
.io_parallelOut_388(dataOut[388]),
.io_parallelOut_389(dataOut[389]),
.io_parallelOut_390(dataOut[390]),
.io_parallelOut_391(dataOut[391]),
.io_parallelOut_392(dataOut[392]),
.io_parallelOut_393(dataOut[393]),
.io_parallelOut_394(dataOut[394]),
.io_parallelOut_395(dataOut[395]),
.io_parallelOut_396(dataOut[396]),
.io_parallelOut_397(dataOut[397]),
.io_parallelOut_398(dataOut[398]),
.io_parallelOut_399(dataOut[399]),
.io_parallelOut_400(dataOut[400]),
.io_parallelOut_401(dataOut[401]),
.io_parallelOut_402(dataOut[402]),
.io_parallelOut_403(dataOut[403]),
.io_parallelOut_404(dataOut[404]),
.io_parallelOut_405(dataOut[405]),
.io_parallelOut_406(dataOut[406]),
.io_parallelOut_407(dataOut[407]),
.io_parallelOut_408(dataOut[408]),
.io_parallelOut_409(dataOut[409]),
.io_parallelOut_410(dataOut[410]),
.io_parallelOut_411(dataOut[411]),
.io_parallelOut_412(dataOut[412]),
.io_parallelOut_413(dataOut[413]),
.io_parallelOut_414(dataOut[414]),
.io_parallelOut_415(dataOut[415]),
.io_parallelOut_416(dataOut[416]),
.io_parallelOut_417(dataOut[417]),
.io_parallelOut_418(dataOut[418]),
.io_parallelOut_419(dataOut[419]),
.io_parallelOut_420(dataOut[420]),
.io_parallelOut_421(dataOut[421]),
.io_parallelOut_422(dataOut[422]),
.io_parallelOut_423(dataOut[423]),
.io_parallelOut_424(dataOut[424]),
.io_parallelOut_425(dataOut[425]),
.io_parallelOut_426(dataOut[426]),
.io_parallelOut_427(dataOut[427]),
.io_parallelOut_428(dataOut[428]),
.io_parallelOut_429(dataOut[429]),
.io_parallelOut_430(dataOut[430]),
.io_parallelOut_431(dataOut[431]),
.io_parallelOut_432(dataOut[432]),
.io_parallelOut_433(dataOut[433]),
.io_parallelOut_434(dataOut[434]),
.io_parallelOut_435(dataOut[435]),
.io_parallelOut_436(dataOut[436]),
.io_parallelOut_437(dataOut[437]),
.io_parallelOut_438(dataOut[438]),
.io_parallelOut_439(dataOut[439]),
.io_parallelOut_440(dataOut[440]),
.io_parallelOut_441(dataOut[441]),
.io_parallelOut_442(dataOut[442]),
.io_parallelOut_443(dataOut[443]),
.io_parallelOut_444(dataOut[444]),
.io_parallelOut_445(dataOut[445]),
.io_parallelOut_446(dataOut[446]),
.io_parallelOut_447(dataOut[447]),
.io_parallelOut_448(dataOut[448]),
.io_parallelOut_449(dataOut[449]),
.io_parallelOut_450(dataOut[450]),
.io_parallelOut_451(dataOut[451]),
.io_parallelOut_452(dataOut[452]),
.io_parallelOut_453(dataOut[453]),
.io_parallelOut_454(dataOut[454]),
.io_parallelOut_455(dataOut[455]),
.io_parallelOut_456(dataOut[456]),
.io_parallelOut_457(dataOut[457]),
.io_parallelOut_458(dataOut[458]),
.io_parallelOut_459(dataOut[459]),
.io_parallelOut_460(dataOut[460]),
.io_parallelOut_461(dataOut[461]),
.io_parallelOut_462(dataOut[462]),
.io_parallelOut_463(dataOut[463]),
.io_parallelOut_464(dataOut[464]),
.io_parallelOut_465(dataOut[465]),
.io_parallelOut_466(dataOut[466]),
.io_parallelOut_467(dataOut[467]),
.io_parallelOut_468(dataOut[468]),
.io_parallelOut_469(dataOut[469]),
.io_parallelOut_470(dataOut[470]),
.io_parallelOut_471(dataOut[471]),
.io_parallelOut_472(dataOut[472]),
.io_parallelOut_473(dataOut[473]),
.io_parallelOut_474(dataOut[474]),
.io_parallelOut_475(dataOut[475]),
.io_parallelOut_476(dataOut[476]),
.io_parallelOut_477(dataOut[477]),
.io_parallelOut_478(dataOut[478]),
.io_parallelOut_479(dataOut[479]),
.io_parallelOut_480(dataOut[480]),
.io_parallelOut_481(dataOut[481]),
.io_parallelOut_482(dataOut[482]),
.io_parallelOut_483(dataOut[483]),
.io_parallelOut_484(dataOut[484]),
.io_parallelOut_485(dataOut[485]),
.io_parallelOut_486(dataOut[486]),
.io_parallelOut_487(dataOut[487]),
.io_parallelOut_488(dataOut[488]),
.io_parallelOut_489(dataOut[489]),
.io_parallelOut_490(dataOut[490]),
.io_parallelOut_491(dataOut[491]),
.io_parallelOut_492(dataOut[492]),
.io_parallelOut_493(dataOut[493]),
.io_parallelOut_494(dataOut[494]),
.io_parallelOut_495(dataOut[495]),
.io_parallelOut_496(dataOut[496]),
.io_parallelOut_497(dataOut[497]),
.io_parallelOut_498(dataOut[498]),
.io_parallelOut_499(dataOut[499]),
.io_parallelOut_500(dataOut[500]),
.io_parallelOut_501(dataOut[501]),
.io_parallelOut_502(dataOut[502]),
.io_parallelOut_503(dataOut[503]),
.io_parallelOut_504(dataOut[504]),
.io_parallelOut_505(dataOut[505]),
.io_parallelOut_506(dataOut[506]),
.io_parallelOut_507(dataOut[507]),
.io_parallelOut_508(dataOut[508]),
.io_parallelOut_509(dataOut[509]),
.io_parallelOut_510(dataOut[510]),
.io_parallelOut_511(dataOut[511]),
.io_parallelOut_512(dataOut[512]),
.io_parallelOut_513(dataOut[513]),
.io_parallelOut_514(dataOut[514]),
.io_parallelOut_515(dataOut[515]),
.io_parallelOut_516(dataOut[516]),
.io_parallelOut_517(dataOut[517]),
.io_parallelOut_518(dataOut[518]),
.io_parallelOut_519(dataOut[519]),
.io_parallelOut_520(dataOut[520]),
.io_parallelOut_521(dataOut[521]),
.io_parallelOut_522(dataOut[522]),
.io_parallelOut_523(dataOut[523]),
.io_parallelOut_524(dataOut[524]),
.io_parallelOut_525(dataOut[525]),
.io_parallelOut_526(dataOut[526]),
.io_parallelOut_527(dataOut[527]),
.io_parallelOut_528(dataOut[528]),
.io_parallelOut_529(dataOut[529]),
.io_parallelOut_530(dataOut[530]),
.io_parallelOut_531(dataOut[531]),
.io_parallelOut_532(dataOut[532]),
.io_parallelOut_533(dataOut[533]),
.io_parallelOut_534(dataOut[534]),
.io_parallelOut_535(dataOut[535]),
.io_parallelOut_536(dataOut[536]),
.io_parallelOut_537(dataOut[537]),
.io_parallelOut_538(dataOut[538]),
.io_parallelOut_539(dataOut[539]),
.io_parallelOut_540(dataOut[540]),
.io_parallelOut_541(dataOut[541]),
.io_parallelOut_542(dataOut[542]),
.io_parallelOut_543(dataOut[543]),
.io_parallelOut_544(dataOut[544]),
.io_parallelOut_545(dataOut[545]),
.io_parallelOut_546(dataOut[546]),
.io_parallelOut_547(dataOut[547]),
.io_parallelOut_548(dataOut[548]),
.io_parallelOut_549(dataOut[549]),
.io_parallelOut_550(dataOut[550]),
.io_parallelOut_551(dataOut[551]),
.io_parallelOut_552(dataOut[552]),
.io_parallelOut_553(dataOut[553]),
.io_parallelOut_554(dataOut[554]),
.io_parallelOut_555(dataOut[555]),
.io_parallelOut_556(dataOut[556]),
.io_parallelOut_557(dataOut[557]),
.io_parallelOut_558(dataOut[558]),
.io_parallelOut_559(dataOut[559]),
.io_parallelOut_560(dataOut[560]),
.io_parallelOut_561(dataOut[561]),
.io_parallelOut_562(dataOut[562]),
.io_parallelOut_563(dataOut[563]),
.io_parallelOut_564(dataOut[564]),
.io_parallelOut_565(dataOut[565]),
.io_parallelOut_566(dataOut[566]),
.io_parallelOut_567(dataOut[567]),
.io_parallelOut_568(dataOut[568]),
.io_parallelOut_569(dataOut[569]),
.io_parallelOut_570(dataOut[570]),
.io_parallelOut_571(dataOut[571]),
.io_parallelOut_572(dataOut[572]),
.io_parallelOut_573(dataOut[573]),
.io_parallelOut_574(dataOut[574]),
.io_parallelOut_575(dataOut[575]),
.io_parallelOut_576(dataOut[576]),
.io_parallelOut_577(dataOut[577]),
.io_parallelOut_578(dataOut[578]),
.io_parallelOut_579(dataOut[579]),
.io_parallelOut_580(dataOut[580]),
.io_parallelOut_581(dataOut[581]),
.io_parallelOut_582(dataOut[582]),
.io_parallelOut_583(dataOut[583]),
.io_parallelOut_584(dataOut[584]),
.io_parallelOut_585(dataOut[585]),
.io_parallelOut_586(dataOut[586]),
.io_parallelOut_587(dataOut[587]),
.io_parallelOut_588(dataOut[588]),
.io_parallelOut_589(dataOut[589]),
.io_parallelOut_590(dataOut[590]),
.io_parallelOut_591(dataOut[591]),
.io_parallelOut_592(dataOut[592]),
.io_parallelOut_593(dataOut[593]),
.io_parallelOut_594(dataOut[594]),
.io_parallelOut_595(dataOut[595]),
.io_parallelOut_596(dataOut[596]),
.io_parallelOut_597(dataOut[597]),
.io_parallelOut_598(dataOut[598]),
.io_parallelOut_599(dataOut[599]),
.io_parallelOut_600(dataOut[600]),
.io_parallelOut_601(dataOut[601]),
.io_parallelOut_602(dataOut[602]),
.io_parallelOut_603(dataOut[603]),
.io_parallelOut_604(dataOut[604]),
.io_parallelOut_605(dataOut[605]),
.io_parallelOut_606(dataOut[606]),
.io_parallelOut_607(dataOut[607]),
.io_parallelOut_608(dataOut[608]),
.io_parallelOut_609(dataOut[609]),
.io_parallelOut_610(dataOut[610]),
.io_parallelOut_611(dataOut[611]),
.io_parallelOut_612(dataOut[612]),
.io_parallelOut_613(dataOut[613]),
.io_parallelOut_614(dataOut[614]),
.io_parallelOut_615(dataOut[615]),
.io_parallelOut_616(dataOut[616]),
.io_parallelOut_617(dataOut[617]),
.io_parallelOut_618(dataOut[618]),
.io_parallelOut_619(dataOut[619]),
.io_parallelOut_620(dataOut[620]),
.io_parallelOut_621(dataOut[621]),
.io_parallelOut_622(dataOut[622]),
.io_parallelOut_623(dataOut[623]),
.io_parallelOut_624(dataOut[624]),
.io_parallelOut_625(dataOut[625]),
.io_parallelOut_626(dataOut[626]),
.io_parallelOut_627(dataOut[627]),
.io_parallelOut_628(dataOut[628]),
.io_parallelOut_629(dataOut[629]),
.io_parallelOut_630(dataOut[630]),
.io_parallelOut_631(dataOut[631]),
.io_parallelOut_632(dataOut[632]),
.io_parallelOut_633(dataOut[633]),
.io_parallelOut_634(dataOut[634]),
.io_parallelOut_635(dataOut[635]),
.io_parallelOut_636(dataOut[636]),
.io_parallelOut_637(dataOut[637]),
.io_parallelOut_638(dataOut[638]),
.io_parallelOut_639(dataOut[639]),
.io_parallelOut_640(dataOut[640]),
.io_parallelOut_641(dataOut[641]),
.io_parallelOut_642(dataOut[642]),
.io_parallelOut_643(dataOut[643]),
.io_parallelOut_644(dataOut[644]),
.io_parallelOut_645(dataOut[645]),
.io_parallelOut_646(dataOut[646]),
.io_parallelOut_647(dataOut[647]),
.io_parallelOut_648(dataOut[648]),
.io_parallelOut_649(dataOut[649]),
.io_parallelOut_650(dataOut[650]),
.io_parallelOut_651(dataOut[651]),
.io_parallelOut_652(dataOut[652]),
.io_parallelOut_653(dataOut[653]),
.io_parallelOut_654(dataOut[654]),
.io_parallelOut_655(dataOut[655]),
.io_parallelOut_656(dataOut[656]),
.io_parallelOut_657(dataOut[657]),
.io_parallelOut_658(dataOut[658]),
.io_parallelOut_659(dataOut[659]),
.io_parallelOut_660(dataOut[660]),
.io_parallelOut_661(dataOut[661]),
.io_parallelOut_662(dataOut[662]),
.io_parallelOut_663(dataOut[663]),
.io_parallelOut_664(dataOut[664]),
.io_parallelOut_665(dataOut[665]),
.io_parallelOut_666(dataOut[666]),
.io_parallelOut_667(dataOut[667]),
.io_parallelOut_668(dataOut[668]),
.io_parallelOut_669(dataOut[669]),
.io_parallelOut_670(dataOut[670]),
.io_parallelOut_671(dataOut[671]),
.io_parallelOut_672(dataOut[672]),
.io_parallelOut_673(dataOut[673]),
.io_parallelOut_674(dataOut[674]),
.io_parallelOut_675(dataOut[675]),
.io_parallelOut_676(dataOut[676]),
.io_parallelOut_677(dataOut[677]),
.io_parallelOut_678(dataOut[678]),
.io_parallelOut_679(dataOut[679]),
.io_parallelOut_680(dataOut[680]),
.io_parallelOut_681(dataOut[681]),
.io_parallelOut_682(dataOut[682]),
.io_parallelOut_683(dataOut[683]),
.io_parallelOut_684(dataOut[684]),
.io_parallelOut_685(dataOut[685]),
.io_parallelOut_686(dataOut[686]),
.io_parallelOut_687(dataOut[687]),
.io_parallelOut_688(dataOut[688]),
.io_parallelOut_689(dataOut[689]),
.io_parallelOut_690(dataOut[690]),
.io_parallelOut_691(dataOut[691]),
.io_parallelOut_692(dataOut[692]),
.io_parallelOut_693(dataOut[693]),
.io_parallelOut_694(dataOut[694]),
.io_parallelOut_695(dataOut[695]),
.io_parallelOut_696(dataOut[696]),
.io_parallelOut_697(dataOut[697]),
.io_parallelOut_698(dataOut[698]),
.io_parallelOut_699(dataOut[699]),
.io_parallelOut_700(dataOut[700]),
.io_parallelOut_701(dataOut[701]),
.io_parallelOut_702(dataOut[702]),
.io_parallelOut_703(dataOut[703]),
.io_parallelOut_704(dataOut[704]),
.io_parallelOut_705(dataOut[705]),
.io_parallelOut_706(dataOut[706]),
.io_parallelOut_707(dataOut[707]),
.io_parallelOut_708(dataOut[708]),
.io_parallelOut_709(dataOut[709]),
.io_parallelOut_710(dataOut[710]),
.io_parallelOut_711(dataOut[711]),
.io_parallelOut_712(dataOut[712]),
.io_parallelOut_713(dataOut[713]),
.io_parallelOut_714(dataOut[714]),
.io_parallelOut_715(dataOut[715]),
.io_parallelOut_716(dataOut[716]),
.io_parallelOut_717(dataOut[717]),
.io_parallelOut_718(dataOut[718]),
.io_parallelOut_719(dataOut[719]),
.io_parallelOut_720(dataOut[720]),
.io_parallelOut_721(dataOut[721]),
.io_parallelOut_722(dataOut[722]),
.io_parallelOut_723(dataOut[723]),
.io_parallelOut_724(dataOut[724]),
.io_parallelOut_725(dataOut[725]),
.io_parallelOut_726(dataOut[726]),
.io_parallelOut_727(dataOut[727]),
.io_parallelOut_728(dataOut[728]),
.io_parallelOut_729(dataOut[729]),
.io_parallelOut_730(dataOut[730]),
.io_parallelOut_731(dataOut[731]),
.io_parallelOut_732(dataOut[732]),
.io_parallelOut_733(dataOut[733]),
.io_parallelOut_734(dataOut[734]),
.io_parallelOut_735(dataOut[735]),
.io_parallelOut_736(dataOut[736]),
.io_parallelOut_737(dataOut[737]),
.io_parallelOut_738(dataOut[738]),
.io_parallelOut_739(dataOut[739]),
.io_parallelOut_740(dataOut[740]),
.io_parallelOut_741(dataOut[741]),
.io_parallelOut_742(dataOut[742]),
.io_parallelOut_743(dataOut[743]),
.io_parallelOut_744(dataOut[744]),
.io_parallelOut_745(dataOut[745]),
.io_parallelOut_746(dataOut[746]),
.io_parallelOut_747(dataOut[747]),
.io_parallelOut_748(dataOut[748]),
.io_parallelOut_749(dataOut[749]),
.io_parallelOut_750(dataOut[750]),
.io_parallelOut_751(dataOut[751]),
.io_parallelOut_752(dataOut[752]),
.io_parallelOut_753(dataOut[753]),
.io_parallelOut_754(dataOut[754]),
.io_parallelOut_755(dataOut[755]),
.io_parallelOut_756(dataOut[756]),
.io_parallelOut_757(dataOut[757]),
.io_parallelOut_758(dataOut[758]),
.io_parallelOut_759(dataOut[759]),
.io_parallelOut_760(dataOut[760]),
.io_parallelOut_761(dataOut[761]),
.io_parallelOut_762(dataOut[762]),
.io_parallelOut_763(dataOut[763]),
.io_parallelOut_764(dataOut[764]),
.io_parallelOut_765(dataOut[765]),
.io_parallelOut_766(dataOut[766]),
.io_parallelOut_767(dataOut[767]),
.io_parallelOut_768(dataOut[768]),
.io_parallelOut_769(dataOut[769]),
.io_parallelOut_770(dataOut[770]),
.io_parallelOut_771(dataOut[771]),
.io_parallelOut_772(dataOut[772]),
.io_parallelOut_773(dataOut[773]),
.io_parallelOut_774(dataOut[774]),
.io_parallelOut_775(dataOut[775]),
.io_parallelOut_776(dataOut[776]),
.io_parallelOut_777(dataOut[777]),
.io_parallelOut_778(dataOut[778]),
.io_parallelOut_779(dataOut[779]),
.io_parallelOut_780(dataOut[780]),
.io_parallelOut_781(dataOut[781]),
.io_parallelOut_782(dataOut[782]),
.io_parallelOut_783(dataOut[783]),
.io_parallelOut_784(dataOut[784]),
.io_parallelOut_785(dataOut[785]),
.io_parallelOut_786(dataOut[786]),
.io_parallelOut_787(dataOut[787]),
.io_parallelOut_788(dataOut[788]),
.io_parallelOut_789(dataOut[789]),
.io_parallelOut_790(dataOut[790]),
.io_parallelOut_791(dataOut[791]),
.io_parallelOut_792(dataOut[792]),
.io_parallelOut_793(dataOut[793]),
.io_parallelOut_794(dataOut[794]),
.io_parallelOut_795(dataOut[795]),
.io_parallelOut_796(dataOut[796]),
.io_parallelOut_797(dataOut[797]),
.io_parallelOut_798(dataOut[798]),
.io_parallelOut_799(dataOut[799]),
.io_parallelOut_800(dataOut[800]),
.io_parallelOut_801(dataOut[801]),
.io_parallelOut_802(dataOut[802]),
.io_parallelOut_803(dataOut[803]),
.io_parallelOut_804(dataOut[804]),
.io_parallelOut_805(dataOut[805]),
.io_parallelOut_806(dataOut[806]),
.io_parallelOut_807(dataOut[807]),
.io_parallelOut_808(dataOut[808]),
.io_parallelOut_809(dataOut[809]),
.io_parallelOut_810(dataOut[810]),
.io_parallelOut_811(dataOut[811]),
.io_parallelOut_812(dataOut[812]),
.io_parallelOut_813(dataOut[813]),
.io_parallelOut_814(dataOut[814]),
.io_parallelOut_815(dataOut[815]),
.io_parallelOut_816(dataOut[816]),
.io_parallelOut_817(dataOut[817]),
.io_parallelOut_818(dataOut[818]),
.io_parallelOut_819(dataOut[819]),
.io_parallelOut_820(dataOut[820]),
.io_parallelOut_821(dataOut[821]),
.io_parallelOut_822(dataOut[822]),
.io_parallelOut_823(dataOut[823]),
.io_parallelOut_824(dataOut[824]),
.io_parallelOut_825(dataOut[825]),
.io_parallelOut_826(dataOut[826]),
.io_parallelOut_827(dataOut[827]),
.io_parallelOut_828(dataOut[828]),
.io_parallelOut_829(dataOut[829]),
.io_parallelOut_830(dataOut[830]),
.io_parallelOut_831(dataOut[831]),
.io_parallelOut_832(dataOut[832]),
.io_parallelOut_833(dataOut[833]),
.io_parallelOut_834(dataOut[834]),
.io_parallelOut_835(dataOut[835]),
.io_parallelOut_836(dataOut[836]),
.io_parallelOut_837(dataOut[837]),
.io_parallelOut_838(dataOut[838]),
.io_parallelOut_839(dataOut[839]),
.io_parallelOut_840(dataOut[840]),
.io_parallelOut_841(dataOut[841]),
.io_parallelOut_842(dataOut[842]),
.io_parallelOut_843(dataOut[843]),
.io_parallelOut_844(dataOut[844]),
.io_parallelOut_845(dataOut[845]),
.io_parallelOut_846(dataOut[846]),
.io_parallelOut_847(dataOut[847]),
.io_parallelOut_848(dataOut[848]),
.io_parallelOut_849(dataOut[849]),
.io_parallelOut_850(dataOut[850]),
.io_parallelOut_851(dataOut[851]),
.io_parallelOut_852(dataOut[852]),
.io_parallelOut_853(dataOut[853]),
.io_parallelOut_854(dataOut[854]),
.io_parallelOut_855(dataOut[855]),
.io_parallelOut_856(dataOut[856]),
.io_parallelOut_857(dataOut[857]),
.io_parallelOut_858(dataOut[858]),
.io_parallelOut_859(dataOut[859]),
.io_parallelOut_860(dataOut[860]),
.io_parallelOut_861(dataOut[861]),
.io_parallelOut_862(dataOut[862]),
.io_parallelOut_863(dataOut[863]),
.io_parallelOut_864(dataOut[864]),
.io_parallelOut_865(dataOut[865]),
.io_parallelOut_866(dataOut[866]),
.io_parallelOut_867(dataOut[867]),
.io_parallelOut_868(dataOut[868]),
.io_parallelOut_869(dataOut[869]),
.io_parallelOut_870(dataOut[870]),
.io_parallelOut_871(dataOut[871]),
.io_parallelOut_872(dataOut[872]),
.io_parallelOut_873(dataOut[873]),
.io_parallelOut_874(dataOut[874]),
.io_parallelOut_875(dataOut[875]),
.io_parallelOut_876(dataOut[876]),
.io_parallelOut_877(dataOut[877]),
.io_parallelOut_878(dataOut[878]),
.io_parallelOut_879(dataOut[879]),
.io_parallelOut_880(dataOut[880]),
.io_parallelOut_881(dataOut[881]),
.io_parallelOut_882(dataOut[882]),
.io_parallelOut_883(dataOut[883]),
.io_parallelOut_884(dataOut[884]),
.io_parallelOut_885(dataOut[885]),
.io_parallelOut_886(dataOut[886]),
.io_parallelOut_887(dataOut[887]),
.io_parallelOut_888(dataOut[888]),
.io_parallelOut_889(dataOut[889]),
.io_parallelOut_890(dataOut[890]),
.io_parallelOut_891(dataOut[891]),
.io_parallelOut_892(dataOut[892]),
.io_parallelOut_893(dataOut[893]),
.io_parallelOut_894(dataOut[894]),
.io_parallelOut_895(dataOut[895]),
.io_parallelOut_896(dataOut[896]),
.io_parallelOut_897(dataOut[897]),
.io_parallelOut_898(dataOut[898]),
.io_parallelOut_899(dataOut[899]),
.io_parallelOut_900(dataOut[900]),
.io_parallelOut_901(dataOut[901]),
.io_parallelOut_902(dataOut[902]),
.io_parallelOut_903(dataOut[903]),
.io_parallelOut_904(dataOut[904]),
.io_parallelOut_905(dataOut[905]),
.io_parallelOut_906(dataOut[906]),
.io_parallelOut_907(dataOut[907]),
.io_parallelOut_908(dataOut[908]),
.io_parallelOut_909(dataOut[909]),
.io_parallelOut_910(dataOut[910]),
.io_parallelOut_911(dataOut[911]),
.io_parallelOut_912(dataOut[912]),
.io_parallelOut_913(dataOut[913]),
.io_parallelOut_914(dataOut[914]),
.io_parallelOut_915(dataOut[915]),
.io_parallelOut_916(dataOut[916]),
.io_parallelOut_917(dataOut[917]),
.io_parallelOut_918(dataOut[918]),
.io_parallelOut_919(dataOut[919]),
.io_parallelOut_920(dataOut[920]),
.io_parallelOut_921(dataOut[921]),
.io_parallelOut_922(dataOut[922]),
.io_parallelOut_923(dataOut[923]),
.io_parallelOut_924(dataOut[924]),
.io_parallelOut_925(dataOut[925]),
.io_parallelOut_926(dataOut[926]),
.io_parallelOut_927(dataOut[927]),
.io_parallelOut_928(dataOut[928]),
.io_parallelOut_929(dataOut[929]),
.io_parallelOut_930(dataOut[930]),
.io_parallelOut_931(dataOut[931]),
.io_parallelOut_932(dataOut[932]),
.io_parallelOut_933(dataOut[933]),
.io_parallelOut_934(dataOut[934]),
.io_parallelOut_935(dataOut[935]),
.io_parallelOut_936(dataOut[936]),
.io_parallelOut_937(dataOut[937]),
.io_parallelOut_938(dataOut[938]),
.io_parallelOut_939(dataOut[939]),
.io_parallelOut_940(dataOut[940]),
.io_parallelOut_941(dataOut[941]),
.io_parallelOut_942(dataOut[942]),
.io_parallelOut_943(dataOut[943]),
.io_parallelOut_944(dataOut[944]),
.io_parallelOut_945(dataOut[945]),
.io_parallelOut_946(dataOut[946]),
.io_parallelOut_947(dataOut[947]),
.io_parallelOut_948(dataOut[948]),
.io_parallelOut_949(dataOut[949]),
.io_parallelOut_950(dataOut[950]),
.io_parallelOut_951(dataOut[951]),
.io_parallelOut_952(dataOut[952]),
.io_parallelOut_953(dataOut[953]),
.io_parallelOut_954(dataOut[954]),
.io_parallelOut_955(dataOut[955]),
.io_parallelOut_956(dataOut[956]),
.io_parallelOut_957(dataOut[957]),
.io_parallelOut_958(dataOut[958]),
.io_parallelOut_959(dataOut[959]),
.io_parallelOut_960(dataOut[960]),
.io_parallelOut_961(dataOut[961]),
.io_parallelOut_962(dataOut[962]),
.io_parallelOut_963(dataOut[963]),
.io_parallelOut_964(dataOut[964]),
.io_parallelOut_965(dataOut[965]),
.io_parallelOut_966(dataOut[966]),
.io_parallelOut_967(dataOut[967]),
.io_parallelOut_968(dataOut[968]),
.io_parallelOut_969(dataOut[969]),
.io_parallelOut_970(dataOut[970]),
.io_parallelOut_971(dataOut[971]),
.io_parallelOut_972(dataOut[972]),
.io_parallelOut_973(dataOut[973]),
.io_parallelOut_974(dataOut[974]),
.io_parallelOut_975(dataOut[975]),
.io_parallelOut_976(dataOut[976]),
.io_parallelOut_977(dataOut[977]),
.io_parallelOut_978(dataOut[978]),
.io_parallelOut_979(dataOut[979]),
.io_parallelOut_980(dataOut[980]),
.io_parallelOut_981(dataOut[981]),
.io_parallelOut_982(dataOut[982]),
.io_parallelOut_983(dataOut[983]),
.io_parallelOut_984(dataOut[984]),
.io_parallelOut_985(dataOut[985]),
.io_parallelOut_986(dataOut[986]),
.io_parallelOut_987(dataOut[987]),
.io_parallelOut_988(dataOut[988]),
.io_parallelOut_989(dataOut[989]),
.io_parallelOut_990(dataOut[990]),
.io_parallelOut_991(dataOut[991]),
.io_parallelOut_992(dataOut[992]),
.io_parallelOut_993(dataOut[993]),
.io_parallelOut_994(dataOut[994]),
.io_parallelOut_995(dataOut[995]),
.io_parallelOut_996(dataOut[996]),
.io_parallelOut_997(dataOut[997]),
.io_parallelOut_998(dataOut[998]),
.io_parallelOut_999(dataOut[999]),
.io_parallelOut_1000(dataOut[1000]),
.io_parallelOut_1001(dataOut[1001]),
.io_parallelOut_1002(dataOut[1002]),
.io_parallelOut_1003(dataOut[1003]),
.io_parallelOut_1004(dataOut[1004]),
.io_parallelOut_1005(dataOut[1005]),
.io_parallelOut_1006(dataOut[1006]),
.io_parallelOut_1007(dataOut[1007]),
.io_parallelOut_1008(dataOut[1008]),
.io_parallelOut_1009(dataOut[1009]),
.io_parallelOut_1010(dataOut[1010]),
.io_parallelOut_1011(dataOut[1011]),
.io_parallelOut_1012(dataOut[1012]),
.io_parallelOut_1013(dataOut[1013]),
.io_parallelOut_1014(dataOut[1014]),
.io_parallelOut_1015(dataOut[1015]),
.io_parallelOut_1016(dataOut[1016]),
.io_parallelOut_1017(dataOut[1017]),
.io_parallelOut_1018(dataOut[1018]),
.io_parallelOut_1019(dataOut[1019]),
.io_parallelOut_1020(dataOut[1020]),
.io_parallelOut_1021(dataOut[1021]),
.io_parallelOut_1022(dataOut[1022]),
.io_parallelOut_1023(dataOut[1023]),
.io_parallelOut_1024(dataOut[1024]),
.io_parallelOut_1025(dataOut[1025]),
.io_parallelOut_1026(dataOut[1026]),
.io_parallelOut_1027(dataOut[1027]),
.io_parallelOut_1028(dataOut[1028]),
.io_parallelOut_1029(dataOut[1029]),
.io_parallelOut_1030(dataOut[1030]),
.io_parallelOut_1031(dataOut[1031]),
.io_parallelOut_1032(dataOut[1032]),
.io_parallelOut_1033(dataOut[1033]),
.io_parallelOut_1034(dataOut[1034]),
.io_parallelOut_1035(dataOut[1035]),
.io_parallelOut_1036(dataOut[1036]),
.io_parallelOut_1037(dataOut[1037]),
.io_parallelOut_1038(dataOut[1038]),
.io_parallelOut_1039(dataOut[1039]),
.io_parallelOut_1040(dataOut[1040]),
.io_parallelOut_1041(dataOut[1041]),
.io_parallelOut_1042(dataOut[1042]),
.io_parallelOut_1043(dataOut[1043]),
.io_parallelOut_1044(dataOut[1044]),
.io_parallelOut_1045(dataOut[1045]),
.io_parallelOut_1046(dataOut[1046]),
.io_parallelOut_1047(dataOut[1047]),
.io_parallelOut_1048(dataOut[1048]),
.io_parallelOut_1049(dataOut[1049]),
.io_parallelOut_1050(dataOut[1050]),
.io_parallelOut_1051(dataOut[1051]),
.io_parallelOut_1052(dataOut[1052]),
.io_parallelOut_1053(dataOut[1053]),
.io_parallelOut_1054(dataOut[1054]),
.io_parallelOut_1055(dataOut[1055]),
.io_parallelOut_1056(dataOut[1056]),
.io_parallelOut_1057(dataOut[1057]),
.io_parallelOut_1058(dataOut[1058]),
.io_parallelOut_1059(dataOut[1059]),
.io_parallelOut_1060(dataOut[1060]),
.io_parallelOut_1061(dataOut[1061]),
.io_parallelOut_1062(dataOut[1062]),
.io_parallelOut_1063(dataOut[1063]),
.io_parallelOut_1064(dataOut[1064]),
.io_parallelOut_1065(dataOut[1065]),
.io_parallelOut_1066(dataOut[1066]),
.io_parallelOut_1067(dataOut[1067]),
.io_parallelOut_1068(dataOut[1068]),
.io_parallelOut_1069(dataOut[1069]),
.io_parallelOut_1070(dataOut[1070]),
.io_parallelOut_1071(dataOut[1071]),
.io_parallelOut_1072(dataOut[1072]),
.io_parallelOut_1073(dataOut[1073]),
.io_parallelOut_1074(dataOut[1074]),
.io_parallelOut_1075(dataOut[1075]),
.io_parallelOut_1076(dataOut[1076]),
.io_parallelOut_1077(dataOut[1077]),
.io_parallelOut_1078(dataOut[1078]),
.io_parallelOut_1079(dataOut[1079]),
.io_parallelOut_1080(dataOut[1080]),
.io_parallelOut_1081(dataOut[1081]),
.io_parallelOut_1082(dataOut[1082]),
.io_parallelOut_1083(dataOut[1083]),
.io_parallelOut_1084(dataOut[1084]),
.io_parallelOut_1085(dataOut[1085]),
.io_parallelOut_1086(dataOut[1086]),
.io_parallelOut_1087(dataOut[1087]),
.io_parallelOut_1088(dataOut[1088]),
.io_parallelOut_1089(dataOut[1089]),
.io_parallelOut_1090(dataOut[1090]),
.io_parallelOut_1091(dataOut[1091]),
.io_parallelOut_1092(dataOut[1092]),
.io_parallelOut_1093(dataOut[1093]),
.io_parallelOut_1094(dataOut[1094]),
.io_parallelOut_1095(dataOut[1095]),
.io_parallelOut_1096(dataOut[1096]),
.io_parallelOut_1097(dataOut[1097]),
.io_parallelOut_1098(dataOut[1098]),
.io_parallelOut_1099(dataOut[1099]),
.io_parallelOut_1100(dataOut[1100]),
.io_parallelOut_1101(dataOut[1101]),
.io_parallelOut_1102(dataOut[1102]),
.io_parallelOut_1103(dataOut[1103]),
.io_parallelOut_1104(dataOut[1104]),
.io_parallelOut_1105(dataOut[1105]),
.io_parallelOut_1106(dataOut[1106]),
.io_parallelOut_1107(dataOut[1107]),
.io_parallelOut_1108(dataOut[1108]),
.io_parallelOut_1109(dataOut[1109]),
.io_parallelOut_1110(dataOut[1110]),
.io_parallelOut_1111(dataOut[1111]),
.io_parallelOut_1112(dataOut[1112]),
.io_parallelOut_1113(dataOut[1113]),
.io_parallelOut_1114(dataOut[1114]),
.io_parallelOut_1115(dataOut[1115]),
.io_parallelOut_1116(dataOut[1116]),
.io_parallelOut_1117(dataOut[1117]),
.io_parallelOut_1118(dataOut[1118]),
.io_parallelOut_1119(dataOut[1119]),
.io_parallelOut_1120(dataOut[1120]),
.io_parallelOut_1121(dataOut[1121]),
.io_parallelOut_1122(dataOut[1122]),
.io_parallelOut_1123(dataOut[1123]),
.io_parallelOut_1124(dataOut[1124]),
.io_parallelOut_1125(dataOut[1125]),
.io_parallelOut_1126(dataOut[1126]),
.io_parallelOut_1127(dataOut[1127]),
.io_parallelOut_1128(dataOut[1128]),
.io_parallelOut_1129(dataOut[1129]),
.io_parallelOut_1130(dataOut[1130]),
.io_parallelOut_1131(dataOut[1131]),
.io_parallelOut_1132(dataOut[1132]),
.io_parallelOut_1133(dataOut[1133]),
.io_parallelOut_1134(dataOut[1134]),
.io_parallelOut_1135(dataOut[1135]),
.io_parallelOut_1136(dataOut[1136]),
.io_parallelOut_1137(dataOut[1137]),
.io_parallelOut_1138(dataOut[1138]),
.io_parallelOut_1139(dataOut[1139]),
.io_parallelOut_1140(dataOut[1140]),
.io_parallelOut_1141(dataOut[1141]),
.io_parallelOut_1142(dataOut[1142]),
.io_parallelOut_1143(dataOut[1143]),
.io_parallelOut_1144(dataOut[1144]),
.io_parallelOut_1145(dataOut[1145]),
.io_parallelOut_1146(dataOut[1146]),
.io_parallelOut_1147(dataOut[1147]),
.io_parallelOut_1148(dataOut[1148]),
.io_parallelOut_1149(dataOut[1149]),
.io_parallelOut_1150(dataOut[1150]),
.io_parallelOut_1151(dataOut[1151]),
.io_parallelOut_1152(dataOut[1152]),
.io_parallelOut_1153(dataOut[1153]),
.io_parallelOut_1154(dataOut[1154]),
.io_parallelOut_1155(dataOut[1155]),
.io_parallelOut_1156(dataOut[1156]),
.io_parallelOut_1157(dataOut[1157]),
.io_parallelOut_1158(dataOut[1158]),
.io_parallelOut_1159(dataOut[1159]),
.io_parallelOut_1160(dataOut[1160]),
.io_parallelOut_1161(dataOut[1161]),
.io_parallelOut_1162(dataOut[1162]),
.io_parallelOut_1163(dataOut[1163]),
.io_parallelOut_1164(dataOut[1164]),
.io_parallelOut_1165(dataOut[1165]),
.io_parallelOut_1166(dataOut[1166]),
.io_parallelOut_1167(dataOut[1167]),
.io_parallelOut_1168(dataOut[1168]),
.io_parallelOut_1169(dataOut[1169]),
.io_parallelOut_1170(dataOut[1170]),
.io_parallelOut_1171(dataOut[1171]),
.io_parallelOut_1172(dataOut[1172]),
.io_parallelOut_1173(dataOut[1173]),
.io_parallelOut_1174(dataOut[1174]),
.io_parallelOut_1175(dataOut[1175]),
.io_parallelOut_1176(dataOut[1176]),
.io_parallelOut_1177(dataOut[1177]),
.io_parallelOut_1178(dataOut[1178]),
.io_parallelOut_1179(dataOut[1179]),
.io_parallelOut_1180(dataOut[1180]),
.io_parallelOut_1181(dataOut[1181]),
.io_parallelOut_1182(dataOut[1182]),
.io_parallelOut_1183(dataOut[1183]),
.io_parallelOut_1184(dataOut[1184]),
.io_parallelOut_1185(dataOut[1185]),
.io_parallelOut_1186(dataOut[1186]),
.io_parallelOut_1187(dataOut[1187]),
.io_parallelOut_1188(dataOut[1188]),
.io_parallelOut_1189(dataOut[1189]),
.io_parallelOut_1190(dataOut[1190]),
.io_parallelOut_1191(dataOut[1191]),
.io_parallelOut_1192(dataOut[1192]),
.io_parallelOut_1193(dataOut[1193]),
.io_parallelOut_1194(dataOut[1194]),
.io_parallelOut_1195(dataOut[1195]),
.io_parallelOut_1196(dataOut[1196]),
.io_parallelOut_1197(dataOut[1197]),
.io_parallelOut_1198(dataOut[1198]),
.io_parallelOut_1199(dataOut[1199]),
.io_parallelOut_1200(dataOut[1200]),
.io_parallelOut_1201(dataOut[1201]),
.io_parallelOut_1202(dataOut[1202]),
.io_parallelOut_1203(dataOut[1203]),
.io_parallelOut_1204(dataOut[1204]),
.io_parallelOut_1205(dataOut[1205]),
.io_parallelOut_1206(dataOut[1206]),
.io_parallelOut_1207(dataOut[1207]),
.io_parallelOut_1208(dataOut[1208]),
.io_parallelOut_1209(dataOut[1209]),
.io_parallelOut_1210(dataOut[1210]),
.io_parallelOut_1211(dataOut[1211]),
.io_parallelOut_1212(dataOut[1212]),
.io_parallelOut_1213(dataOut[1213]),
.io_parallelOut_1214(dataOut[1214]),
.io_parallelOut_1215(dataOut[1215]),
.io_parallelOut_1216(dataOut[1216]),
.io_parallelOut_1217(dataOut[1217]),
.io_parallelOut_1218(dataOut[1218]),
.io_parallelOut_1219(dataOut[1219]),
.io_parallelOut_1220(dataOut[1220]),
.io_parallelOut_1221(dataOut[1221]),
.io_parallelOut_1222(dataOut[1222]),
.io_parallelOut_1223(dataOut[1223]),
.io_parallelOut_1224(dataOut[1224]),
.io_parallelOut_1225(dataOut[1225]),
.io_parallelOut_1226(dataOut[1226]),
.io_parallelOut_1227(dataOut[1227]),
.io_parallelOut_1228(dataOut[1228]),
.io_parallelOut_1229(dataOut[1229]),
.io_parallelOut_1230(dataOut[1230]),
.io_parallelOut_1231(dataOut[1231]),
.io_parallelOut_1232(dataOut[1232]),
.io_parallelOut_1233(dataOut[1233]),
.io_parallelOut_1234(dataOut[1234]),
.io_parallelOut_1235(dataOut[1235]),
.io_parallelOut_1236(dataOut[1236]),
.io_parallelOut_1237(dataOut[1237]),
.io_parallelOut_1238(dataOut[1238]),
.io_parallelOut_1239(dataOut[1239]),
.io_parallelOut_1240(dataOut[1240]),
.io_parallelOut_1241(dataOut[1241]),
.io_parallelOut_1242(dataOut[1242]),
.io_parallelOut_1243(dataOut[1243]),
.io_parallelOut_1244(dataOut[1244]),
.io_parallelOut_1245(dataOut[1245]),
.io_parallelOut_1246(dataOut[1246]),
.io_parallelOut_1247(dataOut[1247]),
.io_parallelOut_1248(dataOut[1248]),
.io_parallelOut_1249(dataOut[1249]),
.io_parallelOut_1250(dataOut[1250]),
.io_parallelOut_1251(dataOut[1251]),
.io_parallelOut_1252(dataOut[1252]),
.io_parallelOut_1253(dataOut[1253]),
.io_parallelOut_1254(dataOut[1254]),
.io_parallelOut_1255(dataOut[1255]),
.io_parallelOut_1256(dataOut[1256]),
.io_parallelOut_1257(dataOut[1257]),
.io_parallelOut_1258(dataOut[1258]),
.io_parallelOut_1259(dataOut[1259]),
.io_parallelOut_1260(dataOut[1260]),
.io_parallelOut_1261(dataOut[1261]),
.io_parallelOut_1262(dataOut[1262]),
.io_parallelOut_1263(dataOut[1263]),
.io_parallelOut_1264(dataOut[1264]),
.io_parallelOut_1265(dataOut[1265]),
.io_parallelOut_1266(dataOut[1266]),
.io_parallelOut_1267(dataOut[1267]),
.io_parallelOut_1268(dataOut[1268]),
.io_parallelOut_1269(dataOut[1269]),
.io_parallelOut_1270(dataOut[1270]),
.io_parallelOut_1271(dataOut[1271]),
.io_parallelOut_1272(dataOut[1272]),
.io_parallelOut_1273(dataOut[1273]),
.io_parallelOut_1274(dataOut[1274]),
.io_parallelOut_1275(dataOut[1275]),
.io_parallelOut_1276(dataOut[1276]),
.io_parallelOut_1277(dataOut[1277]),
.io_parallelOut_1278(dataOut[1278]),
.io_parallelOut_1279(dataOut[1279]),
.io_parallelOut_1280(dataOut[1280]),
.io_parallelOut_1281(dataOut[1281]),
.io_parallelOut_1282(dataOut[1282]),
.io_parallelOut_1283(dataOut[1283]),
.io_parallelOut_1284(dataOut[1284]),
.io_parallelOut_1285(dataOut[1285]),
.io_parallelOut_1286(dataOut[1286]),
.io_parallelOut_1287(dataOut[1287]),
.io_parallelOut_1288(dataOut[1288]),
.io_parallelOut_1289(dataOut[1289]),
.io_parallelOut_1290(dataOut[1290]),
.io_parallelOut_1291(dataOut[1291]),
.io_parallelOut_1292(dataOut[1292]),
.io_parallelOut_1293(dataOut[1293]),
.io_parallelOut_1294(dataOut[1294]),
.io_parallelOut_1295(dataOut[1295]),
.io_parallelOut_1296(dataOut[1296]),
.io_parallelOut_1297(dataOut[1297]),
.io_parallelOut_1298(dataOut[1298]),
.io_parallelOut_1299(dataOut[1299]),
.io_parallelOut_1300(dataOut[1300]),
.io_parallelOut_1301(dataOut[1301]),
.io_parallelOut_1302(dataOut[1302]),
.io_parallelOut_1303(dataOut[1303]),
.io_parallelOut_1304(dataOut[1304]),
.io_parallelOut_1305(dataOut[1305]),
.io_parallelOut_1306(dataOut[1306]),
.io_parallelOut_1307(dataOut[1307]),
.io_parallelOut_1308(dataOut[1308]),
.io_parallelOut_1309(dataOut[1309]),
.io_parallelOut_1310(dataOut[1310]),
.io_parallelOut_1311(dataOut[1311]),
.io_parallelOut_1312(dataOut[1312]),
.io_parallelOut_1313(dataOut[1313]),
.io_parallelOut_1314(dataOut[1314]),
.io_parallelOut_1315(dataOut[1315]),
.io_parallelOut_1316(dataOut[1316]),
.io_parallelOut_1317(dataOut[1317]),
.io_parallelOut_1318(dataOut[1318]),
.io_parallelOut_1319(dataOut[1319]),
.io_parallelOut_1320(dataOut[1320]),
.io_parallelOut_1321(dataOut[1321]),
.io_parallelOut_1322(dataOut[1322]),
.io_parallelOut_1323(dataOut[1323]),
.io_parallelOut_1324(dataOut[1324]),
.io_parallelOut_1325(dataOut[1325]),
.io_parallelOut_1326(dataOut[1326]),
.io_parallelOut_1327(dataOut[1327]),
.io_parallelOut_1328(dataOut[1328]),
.io_parallelOut_1329(dataOut[1329]),
.io_parallelOut_1330(dataOut[1330]),
.io_parallelOut_1331(dataOut[1331]),
.io_parallelOut_1332(dataOut[1332]),
.io_parallelOut_1333(dataOut[1333]),
.io_parallelOut_1334(dataOut[1334]),
.io_parallelOut_1335(dataOut[1335]),
.io_parallelOut_1336(dataOut[1336]),
.io_parallelOut_1337(dataOut[1337]),
.io_parallelOut_1338(dataOut[1338]),
.io_parallelOut_1339(dataOut[1339]),
.io_parallelOut_1340(dataOut[1340]),
.io_parallelOut_1341(dataOut[1341]),
.io_parallelOut_1342(dataOut[1342]),
.io_parallelOut_1343(dataOut[1343]),
.io_parallelOut_1344(dataOut[1344]),
.io_parallelOut_1345(dataOut[1345]),
.io_parallelOut_1346(dataOut[1346]),
.io_parallelOut_1347(dataOut[1347]),
.io_parallelOut_1348(dataOut[1348]),
.io_parallelOut_1349(dataOut[1349]),
.io_parallelOut_1350(dataOut[1350]),
.io_parallelOut_1351(dataOut[1351]),
.io_parallelOut_1352(dataOut[1352]),
.io_parallelOut_1353(dataOut[1353]),
.io_parallelOut_1354(dataOut[1354]),
.io_parallelOut_1355(dataOut[1355]),
.io_parallelOut_1356(dataOut[1356]),
.io_parallelOut_1357(dataOut[1357]),
.io_parallelOut_1358(dataOut[1358]),
.io_parallelOut_1359(dataOut[1359]),
.io_parallelOut_1360(dataOut[1360]),
.io_parallelOut_1361(dataOut[1361]),
.io_parallelOut_1362(dataOut[1362]),
.io_parallelOut_1363(dataOut[1363]),
.io_parallelOut_1364(dataOut[1364]),
.io_parallelOut_1365(dataOut[1365]),
.io_parallelOut_1366(dataOut[1366]),
.io_parallelOut_1367(dataOut[1367]),
.io_parallelOut_1368(dataOut[1368]),
.io_parallelOut_1369(dataOut[1369]),
.io_parallelOut_1370(dataOut[1370]),
.io_parallelOut_1371(dataOut[1371]),
.io_parallelOut_1372(dataOut[1372]),
.io_parallelOut_1373(dataOut[1373]),
.io_parallelOut_1374(dataOut[1374]),
.io_parallelOut_1375(dataOut[1375]),
.io_parallelOut_1376(dataOut[1376]),
.io_parallelOut_1377(dataOut[1377]),
.io_parallelOut_1378(dataOut[1378]),
.io_parallelOut_1379(dataOut[1379]),
.io_parallelOut_1380(dataOut[1380]),
.io_parallelOut_1381(dataOut[1381]),
.io_parallelOut_1382(dataOut[1382]),
.io_parallelOut_1383(dataOut[1383]),
.io_parallelOut_1384(dataOut[1384]),
.io_parallelOut_1385(dataOut[1385]),
.io_parallelOut_1386(dataOut[1386]),
.io_parallelOut_1387(dataOut[1387]),
.io_parallelOut_1388(dataOut[1388]),
.io_parallelOut_1389(dataOut[1389]),
.io_parallelOut_1390(dataOut[1390]),
.io_parallelOut_1391(dataOut[1391]),
.io_parallelOut_1392(dataOut[1392]),
.io_parallelOut_1393(dataOut[1393]),
.io_parallelOut_1394(dataOut[1394]),
.io_parallelOut_1395(dataOut[1395]),
.io_parallelOut_1396(dataOut[1396]),
.io_parallelOut_1397(dataOut[1397]),
.io_parallelOut_1398(dataOut[1398]),
.io_parallelOut_1399(dataOut[1399]),
.io_parallelOut_1400(dataOut[1400]),
.io_parallelOut_1401(dataOut[1401]),
.io_parallelOut_1402(dataOut[1402]),
.io_parallelOut_1403(dataOut[1403]),
.io_parallelOut_1404(dataOut[1404]),
.io_parallelOut_1405(dataOut[1405]),
.io_parallelOut_1406(dataOut[1406]),
.io_parallelOut_1407(dataOut[1407]),
.io_parallelOut_1408(dataOut[1408]),
.io_parallelOut_1409(dataOut[1409]),
.io_parallelOut_1410(dataOut[1410]),
.io_parallelOut_1411(dataOut[1411]),
.io_parallelOut_1412(dataOut[1412]),
.io_parallelOut_1413(dataOut[1413]),
.io_parallelOut_1414(dataOut[1414]),
.io_parallelOut_1415(dataOut[1415]),
.io_parallelOut_1416(dataOut[1416]),
.io_parallelOut_1417(dataOut[1417]),
.io_parallelOut_1418(dataOut[1418]),
.io_parallelOut_1419(dataOut[1419]),
.io_parallelOut_1420(dataOut[1420]),
.io_parallelOut_1421(dataOut[1421]),
.io_parallelOut_1422(dataOut[1422]),
.io_parallelOut_1423(dataOut[1423]),
.io_parallelOut_1424(dataOut[1424]),
.io_parallelOut_1425(dataOut[1425]),
.io_parallelOut_1426(dataOut[1426]),
.io_parallelOut_1427(dataOut[1427]),
.io_parallelOut_1428(dataOut[1428]),
.io_parallelOut_1429(dataOut[1429]),
.io_parallelOut_1430(dataOut[1430]),
.io_parallelOut_1431(dataOut[1431]),
.io_parallelOut_1432(dataOut[1432]),
.io_parallelOut_1433(dataOut[1433]),
.io_parallelOut_1434(dataOut[1434]),
.io_parallelOut_1435(dataOut[1435]),
.io_parallelOut_1436(dataOut[1436]),
.io_parallelOut_1437(dataOut[1437]),
.io_parallelOut_1438(dataOut[1438]),
.io_parallelOut_1439(dataOut[1439]),
.io_parallelOut_1440(dataOut[1440]),
.io_parallelOut_1441(dataOut[1441]),
.io_parallelOut_1442(dataOut[1442]),
.io_parallelOut_1443(dataOut[1443]),
.io_parallelOut_1444(dataOut[1444]),
.io_parallelOut_1445(dataOut[1445]),
.io_parallelOut_1446(dataOut[1446]),
.io_parallelOut_1447(dataOut[1447]),
.io_parallelOut_1448(dataOut[1448]),
.io_parallelOut_1449(dataOut[1449]),
.io_parallelOut_1450(dataOut[1450]),
.io_parallelOut_1451(dataOut[1451]),
.io_parallelOut_1452(dataOut[1452]),
.io_parallelOut_1453(dataOut[1453]),
.io_parallelOut_1454(dataOut[1454]),
.io_parallelOut_1455(dataOut[1455]),
.io_parallelOut_1456(dataOut[1456]),
.io_parallelOut_1457(dataOut[1457]),
.io_parallelOut_1458(dataOut[1458]),
.io_parallelOut_1459(dataOut[1459]),
.io_parallelOut_1460(dataOut[1460]),
.io_parallelOut_1461(dataOut[1461]),
.io_parallelOut_1462(dataOut[1462]),
.io_parallelOut_1463(dataOut[1463]),
.io_parallelOut_1464(dataOut[1464]),
.io_parallelOut_1465(dataOut[1465]),
.io_parallelOut_1466(dataOut[1466]),
.io_parallelOut_1467(dataOut[1467]),
.io_parallelOut_1468(dataOut[1468]),
.io_parallelOut_1469(dataOut[1469]),
.io_parallelOut_1470(dataOut[1470]),
.io_parallelOut_1471(dataOut[1471]),
.io_parallelOut_1472(dataOut[1472]),
.io_parallelOut_1473(dataOut[1473]),
.io_parallelOut_1474(dataOut[1474]),
.io_parallelOut_1475(dataOut[1475]),
.io_parallelOut_1476(dataOut[1476]),
.io_parallelOut_1477(dataOut[1477]),
.io_parallelOut_1478(dataOut[1478]),
.io_parallelOut_1479(dataOut[1479]),
.io_parallelOut_1480(dataOut[1480]),
.io_parallelOut_1481(dataOut[1481]),
.io_parallelOut_1482(dataOut[1482]),
.io_parallelOut_1483(dataOut[1483]),
.io_parallelOut_1484(dataOut[1484]),
.io_parallelOut_1485(dataOut[1485]),
.io_parallelOut_1486(dataOut[1486]),
.io_parallelOut_1487(dataOut[1487]),
.io_parallelOut_1488(dataOut[1488]),
.io_parallelOut_1489(dataOut[1489]),
.io_parallelOut_1490(dataOut[1490]),
.io_parallelOut_1491(dataOut[1491]),
.io_parallelOut_1492(dataOut[1492]),
.io_parallelOut_1493(dataOut[1493]),
.io_parallelOut_1494(dataOut[1494]),
.io_parallelOut_1495(dataOut[1495]),
.io_parallelOut_1496(dataOut[1496]),
.io_parallelOut_1497(dataOut[1497]),
.io_parallelOut_1498(dataOut[1498]),
.io_parallelOut_1499(dataOut[1499]),
.io_parallelOut_1500(dataOut[1500]),
.io_parallelOut_1501(dataOut[1501]),
.io_parallelOut_1502(dataOut[1502]),
.io_parallelOut_1503(dataOut[1503]),
.io_parallelOut_1504(dataOut[1504]),
.io_parallelOut_1505(dataOut[1505]),
.io_parallelOut_1506(dataOut[1506]),
.io_parallelOut_1507(dataOut[1507]),
.io_parallelOut_1508(dataOut[1508]),
.io_parallelOut_1509(dataOut[1509]),
.io_parallelOut_1510(dataOut[1510]),
.io_parallelOut_1511(dataOut[1511]),
.io_parallelOut_1512(dataOut[1512]),
.io_parallelOut_1513(dataOut[1513]),
.io_parallelOut_1514(dataOut[1514]),
.io_parallelOut_1515(dataOut[1515]),
.io_parallelOut_1516(dataOut[1516]),
.io_parallelOut_1517(dataOut[1517]),
.io_parallelOut_1518(dataOut[1518]),
.io_parallelOut_1519(dataOut[1519]),
.io_parallelOut_1520(dataOut[1520]),
.io_parallelOut_1521(dataOut[1521]),
.io_parallelOut_1522(dataOut[1522]),
.io_parallelOut_1523(dataOut[1523]),
.io_parallelOut_1524(dataOut[1524]),
.io_parallelOut_1525(dataOut[1525]),
.io_parallelOut_1526(dataOut[1526]),
.io_parallelOut_1527(dataOut[1527]),
.io_parallelOut_1528(dataOut[1528]),
.io_parallelOut_1529(dataOut[1529]),
.io_parallelOut_1530(dataOut[1530]),
.io_parallelOut_1531(dataOut[1531]),
.io_parallelOut_1532(dataOut[1532]),
.io_parallelOut_1533(dataOut[1533]),
.io_parallelOut_1534(dataOut[1534]),
.io_parallelOut_1535(dataOut[1535]),
.io_parallelOut_1536(dataOut[1536]),
.io_parallelOut_1537(dataOut[1537]),
.io_parallelOut_1538(dataOut[1538]),
.io_parallelOut_1539(dataOut[1539]),
.io_parallelOut_1540(dataOut[1540]),
.io_parallelOut_1541(dataOut[1541]),
.io_parallelOut_1542(dataOut[1542]),
.io_parallelOut_1543(dataOut[1543]),
.io_parallelOut_1544(dataOut[1544]),
.io_parallelOut_1545(dataOut[1545]),
.io_parallelOut_1546(dataOut[1546]),
.io_parallelOut_1547(dataOut[1547]),
.io_parallelOut_1548(dataOut[1548]),
.io_parallelOut_1549(dataOut[1549]),
.io_parallelOut_1550(dataOut[1550]),
.io_parallelOut_1551(dataOut[1551]),
.io_parallelOut_1552(dataOut[1552]),
.io_parallelOut_1553(dataOut[1553]),
.io_parallelOut_1554(dataOut[1554]),
.io_parallelOut_1555(dataOut[1555]),
.io_parallelOut_1556(dataOut[1556]),
.io_parallelOut_1557(dataOut[1557]),
.io_parallelOut_1558(dataOut[1558]),
.io_parallelOut_1559(dataOut[1559]),
.io_parallelOut_1560(dataOut[1560]),
.io_parallelOut_1561(dataOut[1561]),
.io_parallelOut_1562(dataOut[1562]),
.io_parallelOut_1563(dataOut[1563]),
.io_parallelOut_1564(dataOut[1564]),
.io_parallelOut_1565(dataOut[1565]),
.io_parallelOut_1566(dataOut[1566]),
.io_parallelOut_1567(dataOut[1567]),
.io_parallelOut_1568(dataOut[1568]),
.io_parallelOut_1569(dataOut[1569]),
.io_parallelOut_1570(dataOut[1570]),
.io_parallelOut_1571(dataOut[1571]),
.io_parallelOut_1572(dataOut[1572]),
.io_parallelOut_1573(dataOut[1573]),
.io_parallelOut_1574(dataOut[1574]),
.io_parallelOut_1575(dataOut[1575]),
.io_parallelOut_1576(dataOut[1576]),
.io_parallelOut_1577(dataOut[1577]),
.io_parallelOut_1578(dataOut[1578]),
.io_parallelOut_1579(dataOut[1579]),
.io_parallelOut_1580(dataOut[1580]),
.io_parallelOut_1581(dataOut[1581]),
.io_parallelOut_1582(dataOut[1582]),
.io_parallelOut_1583(dataOut[1583]),
.io_parallelOut_1584(dataOut[1584]),
.io_parallelOut_1585(dataOut[1585]),
.io_parallelOut_1586(dataOut[1586]),
.io_parallelOut_1587(dataOut[1587]),
.io_parallelOut_1588(dataOut[1588]),
.io_parallelOut_1589(dataOut[1589]),
.io_parallelOut_1590(dataOut[1590]),
.io_parallelOut_1591(dataOut[1591]),
.io_parallelOut_1592(dataOut[1592]),
.io_parallelOut_1593(dataOut[1593]),
.io_parallelOut_1594(dataOut[1594]),
.io_parallelOut_1595(dataOut[1595]),
.io_parallelOut_1596(dataOut[1596]),
.io_parallelOut_1597(dataOut[1597]),
.io_parallelOut_1598(dataOut[1598]),
.io_parallelOut_1599(dataOut[1599]),
.io_parallelOut_1600(dataOut[1600]),
.io_parallelOut_1601(dataOut[1601]),
.io_parallelOut_1602(dataOut[1602]),
.io_parallelOut_1603(dataOut[1603]),
.io_parallelOut_1604(dataOut[1604]),
.io_parallelOut_1605(dataOut[1605]),
.io_parallelOut_1606(dataOut[1606]),
.io_parallelOut_1607(dataOut[1607]),
.io_parallelOut_1608(dataOut[1608]),
.io_parallelOut_1609(dataOut[1609]),
.io_parallelOut_1610(dataOut[1610]),
.io_parallelOut_1611(dataOut[1611]),
.io_parallelOut_1612(dataOut[1612]),
.io_parallelOut_1613(dataOut[1613]),
.io_parallelOut_1614(dataOut[1614]),
.io_parallelOut_1615(dataOut[1615]),
.io_parallelOut_1616(dataOut[1616]),
.io_parallelOut_1617(dataOut[1617]),
.io_parallelOut_1618(dataOut[1618]),
.io_parallelOut_1619(dataOut[1619]),
.io_parallelOut_1620(dataOut[1620]),
.io_parallelOut_1621(dataOut[1621]),
.io_parallelOut_1622(dataOut[1622]),
.io_parallelOut_1623(dataOut[1623]),
.io_parallelOut_1624(dataOut[1624]),
.io_parallelOut_1625(dataOut[1625]),
.io_parallelOut_1626(dataOut[1626]),
.io_parallelOut_1627(dataOut[1627]),
.io_parallelOut_1628(dataOut[1628]),
.io_parallelOut_1629(dataOut[1629]),
.io_parallelOut_1630(dataOut[1630]),
.io_parallelOut_1631(dataOut[1631]),
.io_parallelOut_1632(dataOut[1632]),
.io_parallelOut_1633(dataOut[1633]),
.io_parallelOut_1634(dataOut[1634]),
.io_parallelOut_1635(dataOut[1635]),
.io_parallelOut_1636(dataOut[1636]),
.io_parallelOut_1637(dataOut[1637]),
.io_parallelOut_1638(dataOut[1638]),
.io_parallelOut_1639(dataOut[1639]),
.io_parallelOut_1640(dataOut[1640]),
.io_parallelOut_1641(dataOut[1641]),
.io_parallelOut_1642(dataOut[1642]),
.io_parallelOut_1643(dataOut[1643]),
.io_parallelOut_1644(dataOut[1644]),
.io_parallelOut_1645(dataOut[1645]),
.io_parallelOut_1646(dataOut[1646]),
.io_parallelOut_1647(dataOut[1647]),
.io_parallelOut_1648(dataOut[1648]),
.io_parallelOut_1649(dataOut[1649]),
.io_parallelOut_1650(dataOut[1650]),
.io_parallelOut_1651(dataOut[1651]),
.io_parallelOut_1652(dataOut[1652]),
.io_parallelOut_1653(dataOut[1653]),
.io_parallelOut_1654(dataOut[1654]),
.io_parallelOut_1655(dataOut[1655]),
.io_parallelOut_1656(dataOut[1656]),
.io_parallelOut_1657(dataOut[1657]),
.io_parallelOut_1658(dataOut[1658]),
.io_parallelOut_1659(dataOut[1659]),
.io_parallelOut_1660(dataOut[1660]),
.io_parallelOut_1661(dataOut[1661]),
.io_parallelOut_1662(dataOut[1662]),
.io_parallelOut_1663(dataOut[1663]),
.io_parallelOut_1664(dataOut[1664]),
.io_parallelOut_1665(dataOut[1665]),
.io_parallelOut_1666(dataOut[1666]),
.io_parallelOut_1667(dataOut[1667]),
.io_parallelOut_1668(dataOut[1668]),
.io_parallelOut_1669(dataOut[1669]),
.io_parallelOut_1670(dataOut[1670]),
.io_parallelOut_1671(dataOut[1671]),
.io_parallelOut_1672(dataOut[1672]),
.io_parallelOut_1673(dataOut[1673]),
.io_parallelOut_1674(dataOut[1674]),
.io_parallelOut_1675(dataOut[1675]),
.io_parallelOut_1676(dataOut[1676]),
.io_parallelOut_1677(dataOut[1677]),
.io_parallelOut_1678(dataOut[1678]),
.io_parallelOut_1679(dataOut[1679]),
.io_parallelOut_1680(dataOut[1680]),
.io_parallelOut_1681(dataOut[1681]),
.io_parallelOut_1682(dataOut[1682]),
.io_parallelOut_1683(dataOut[1683]),
.io_parallelOut_1684(dataOut[1684]),
.io_parallelOut_1685(dataOut[1685]),
.io_parallelOut_1686(dataOut[1686]),
.io_parallelOut_1687(dataOut[1687]),
.io_parallelOut_1688(dataOut[1688]),
.io_parallelOut_1689(dataOut[1689]),
.io_parallelOut_1690(dataOut[1690]),
.io_parallelOut_1691(dataOut[1691]),
.io_parallelOut_1692(dataOut[1692]),
.io_parallelOut_1693(dataOut[1693]),
.io_parallelOut_1694(dataOut[1694]),
.io_parallelOut_1695(dataOut[1695]),
.io_parallelOut_1696(dataOut[1696]),
.io_parallelOut_1697(dataOut[1697]),
.io_parallelOut_1698(dataOut[1698]),
.io_parallelOut_1699(dataOut[1699]),
.io_parallelOut_1700(dataOut[1700]),
.io_parallelOut_1701(dataOut[1701]),
.io_parallelOut_1702(dataOut[1702]),
.io_parallelOut_1703(dataOut[1703]),
.io_parallelOut_1704(dataOut[1704]),
.io_parallelOut_1705(dataOut[1705]),
.io_parallelOut_1706(dataOut[1706]),
.io_parallelOut_1707(dataOut[1707]),
.io_parallelOut_1708(dataOut[1708]),
.io_parallelOut_1709(dataOut[1709]),
.io_parallelOut_1710(dataOut[1710]),
.io_parallelOut_1711(dataOut[1711]),
.io_parallelOut_1712(dataOut[1712]),
.io_parallelOut_1713(dataOut[1713]),
.io_parallelOut_1714(dataOut[1714]),
.io_parallelOut_1715(dataOut[1715]),
.io_parallelOut_1716(dataOut[1716]),
.io_parallelOut_1717(dataOut[1717]),
.io_parallelOut_1718(dataOut[1718]),
.io_parallelOut_1719(dataOut[1719]),
.io_parallelOut_1720(dataOut[1720]),
.io_parallelOut_1721(dataOut[1721]),
.io_parallelOut_1722(dataOut[1722]),
.io_parallelOut_1723(dataOut[1723]),
.io_parallelOut_1724(dataOut[1724]),
.io_parallelOut_1725(dataOut[1725]),
.io_parallelOut_1726(dataOut[1726]),
.io_parallelOut_1727(dataOut[1727]),
.io_parallelOut_1728(dataOut[1728]),
.io_parallelOut_1729(dataOut[1729]),
.io_parallelOut_1730(dataOut[1730]),
.io_parallelOut_1731(dataOut[1731]),
.io_parallelOut_1732(dataOut[1732]),
.io_parallelOut_1733(dataOut[1733]),
.io_parallelOut_1734(dataOut[1734]),
.io_parallelOut_1735(dataOut[1735]),
.io_parallelOut_1736(dataOut[1736]),
.io_parallelOut_1737(dataOut[1737]),
.io_parallelOut_1738(dataOut[1738]),
.io_parallelOut_1739(dataOut[1739]),
.io_parallelOut_1740(dataOut[1740]),
.io_parallelOut_1741(dataOut[1741]),
.io_parallelOut_1742(dataOut[1742]),
.io_parallelOut_1743(dataOut[1743]),
.io_parallelOut_1744(dataOut[1744]),
.io_parallelOut_1745(dataOut[1745]),
.io_parallelOut_1746(dataOut[1746]),
.io_parallelOut_1747(dataOut[1747]),
.io_parallelOut_1748(dataOut[1748]),
.io_parallelOut_1749(dataOut[1749]),
.io_parallelOut_1750(dataOut[1750]),
.io_parallelOut_1751(dataOut[1751]),
.io_parallelOut_1752(dataOut[1752]),
.io_parallelOut_1753(dataOut[1753]),
.io_parallelOut_1754(dataOut[1754]),
.io_parallelOut_1755(dataOut[1755]),
.io_parallelOut_1756(dataOut[1756]),
.io_parallelOut_1757(dataOut[1757]),
.io_parallelOut_1758(dataOut[1758]),
.io_parallelOut_1759(dataOut[1759]),
.io_parallelOut_1760(dataOut[1760]),
.io_parallelOut_1761(dataOut[1761]),
.io_parallelOut_1762(dataOut[1762]),
.io_parallelOut_1763(dataOut[1763]),
.io_parallelOut_1764(dataOut[1764]),
.io_parallelOut_1765(dataOut[1765]),
.io_parallelOut_1766(dataOut[1766]),
.io_parallelOut_1767(dataOut[1767]),
.io_parallelOut_1768(dataOut[1768]),
.io_parallelOut_1769(dataOut[1769]),
.io_parallelOut_1770(dataOut[1770]),
.io_parallelOut_1771(dataOut[1771]),
.io_parallelOut_1772(dataOut[1772]),
.io_parallelOut_1773(dataOut[1773]),
.io_parallelOut_1774(dataOut[1774]),
.io_parallelOut_1775(dataOut[1775]),
.io_parallelOut_1776(dataOut[1776]),
.io_parallelOut_1777(dataOut[1777]),
.io_parallelOut_1778(dataOut[1778]),
.io_parallelOut_1779(dataOut[1779]),
.io_parallelOut_1780(dataOut[1780]),
.io_parallelOut_1781(dataOut[1781]),
.io_parallelOut_1782(dataOut[1782]),
.io_parallelOut_1783(dataOut[1783]),
.io_parallelOut_1784(dataOut[1784]),
.io_parallelOut_1785(dataOut[1785]),
.io_parallelOut_1786(dataOut[1786]),
.io_parallelOut_1787(dataOut[1787]),
.io_parallelOut_1788(dataOut[1788]),
.io_parallelOut_1789(dataOut[1789]),
.io_parallelOut_1790(dataOut[1790]),
.io_parallelOut_1791(dataOut[1791]),
.io_parallelOut_1792(dataOut[1792]),
.io_parallelOut_1793(dataOut[1793]),
.io_parallelOut_1794(dataOut[1794]),
.io_parallelOut_1795(dataOut[1795]),
.io_parallelOut_1796(dataOut[1796]),
.io_parallelOut_1797(dataOut[1797]),
.io_parallelOut_1798(dataOut[1798]),
.io_parallelOut_1799(dataOut[1799]),
.io_parallelOut_1800(dataOut[1800]),
.io_parallelOut_1801(dataOut[1801]),
.io_parallelOut_1802(dataOut[1802]),
.io_parallelOut_1803(dataOut[1803]),
.io_parallelOut_1804(dataOut[1804]),
.io_parallelOut_1805(dataOut[1805]),
.io_parallelOut_1806(dataOut[1806]),
.io_parallelOut_1807(dataOut[1807]),
.io_parallelOut_1808(dataOut[1808]),
.io_parallelOut_1809(dataOut[1809]),
.io_parallelOut_1810(dataOut[1810]),
.io_parallelOut_1811(dataOut[1811]),
.io_parallelOut_1812(dataOut[1812]),
.io_parallelOut_1813(dataOut[1813]),
.io_parallelOut_1814(dataOut[1814]),
.io_parallelOut_1815(dataOut[1815]),
.io_parallelOut_1816(dataOut[1816]),
.io_parallelOut_1817(dataOut[1817]),
.io_parallelOut_1818(dataOut[1818]),
.io_parallelOut_1819(dataOut[1819]),
.io_parallelOut_1820(dataOut[1820]),
.io_parallelOut_1821(dataOut[1821]),
.io_parallelOut_1822(dataOut[1822]),
.io_parallelOut_1823(dataOut[1823]),
.io_parallelOut_1824(dataOut[1824]),
.io_parallelOut_1825(dataOut[1825]),
.io_parallelOut_1826(dataOut[1826]),
.io_parallelOut_1827(dataOut[1827]),
.io_parallelOut_1828(dataOut[1828]),
.io_parallelOut_1829(dataOut[1829]),
.io_parallelOut_1830(dataOut[1830]),
.io_parallelOut_1831(dataOut[1831]),
.io_parallelOut_1832(dataOut[1832]),
.io_parallelOut_1833(dataOut[1833]),
.io_parallelOut_1834(dataOut[1834]),
.io_parallelOut_1835(dataOut[1835]),
.io_parallelOut_1836(dataOut[1836]),
.io_parallelOut_1837(dataOut[1837]),
.io_parallelOut_1838(dataOut[1838]),
.io_parallelOut_1839(dataOut[1839]),
.io_parallelOut_1840(dataOut[1840]),
.io_parallelOut_1841(dataOut[1841]),
.io_parallelOut_1842(dataOut[1842]),
.io_parallelOut_1843(dataOut[1843]),
.io_parallelOut_1844(dataOut[1844]),
.io_parallelOut_1845(dataOut[1845]),
.io_parallelOut_1846(dataOut[1846]),
.io_parallelOut_1847(dataOut[1847]),
.io_parallelOut_1848(dataOut[1848]),
.io_parallelOut_1849(dataOut[1849]),
.io_parallelOut_1850(dataOut[1850]),
.io_parallelOut_1851(dataOut[1851]),
.io_parallelOut_1852(dataOut[1852]),
.io_parallelOut_1853(dataOut[1853]),
.io_parallelOut_1854(dataOut[1854]),
.io_parallelOut_1855(dataOut[1855]),
.io_parallelOut_1856(dataOut[1856]),
.io_parallelOut_1857(dataOut[1857]),
.io_parallelOut_1858(dataOut[1858]),
.io_parallelOut_1859(dataOut[1859]),
.io_parallelOut_1860(dataOut[1860]),
.io_parallelOut_1861(dataOut[1861]),
.io_parallelOut_1862(dataOut[1862]),
.io_parallelOut_1863(dataOut[1863]),
.io_parallelOut_1864(dataOut[1864]),
.io_parallelOut_1865(dataOut[1865]),
.io_parallelOut_1866(dataOut[1866]),
.io_parallelOut_1867(dataOut[1867]),
.io_parallelOut_1868(dataOut[1868]),
.io_parallelOut_1869(dataOut[1869]),
.io_parallelOut_1870(dataOut[1870]),
.io_parallelOut_1871(dataOut[1871]),
.io_parallelOut_1872(dataOut[1872]),
.io_parallelOut_1873(dataOut[1873]),
.io_parallelOut_1874(dataOut[1874]),
.io_parallelOut_1875(dataOut[1875]),
.io_parallelOut_1876(dataOut[1876]),
.io_parallelOut_1877(dataOut[1877]),
.io_parallelOut_1878(dataOut[1878]),
.io_parallelOut_1879(dataOut[1879]),
.io_parallelOut_1880(dataOut[1880]),
.io_parallelOut_1881(dataOut[1881]),
.io_parallelOut_1882(dataOut[1882]),
.io_parallelOut_1883(dataOut[1883]),
.io_parallelOut_1884(dataOut[1884]),
.io_parallelOut_1885(dataOut[1885]),
.io_parallelOut_1886(dataOut[1886]),
.io_parallelOut_1887(dataOut[1887]),
.io_parallelOut_1888(dataOut[1888]),
.io_parallelOut_1889(dataOut[1889]),
.io_parallelOut_1890(dataOut[1890]),
.io_parallelOut_1891(dataOut[1891]),
.io_parallelOut_1892(dataOut[1892]),
.io_parallelOut_1893(dataOut[1893]),
.io_parallelOut_1894(dataOut[1894]),
.io_parallelOut_1895(dataOut[1895]),
.io_parallelOut_1896(dataOut[1896]),
.io_parallelOut_1897(dataOut[1897]),
.io_parallelOut_1898(dataOut[1898]),
.io_parallelOut_1899(dataOut[1899]),
.io_parallelOut_1900(dataOut[1900]),
.io_parallelOut_1901(dataOut[1901]),
.io_parallelOut_1902(dataOut[1902]),
.io_parallelOut_1903(dataOut[1903]),
.io_parallelOut_1904(dataOut[1904]),
.io_parallelOut_1905(dataOut[1905]),
.io_parallelOut_1906(dataOut[1906]),
.io_parallelOut_1907(dataOut[1907]),
.io_parallelOut_1908(dataOut[1908]),
.io_parallelOut_1909(dataOut[1909]),
.io_parallelOut_1910(dataOut[1910]),
.io_parallelOut_1911(dataOut[1911]),
.io_parallelOut_1912(dataOut[1912]),
.io_parallelOut_1913(dataOut[1913]),
.io_parallelOut_1914(dataOut[1914]),
.io_parallelOut_1915(dataOut[1915]),
.io_parallelOut_1916(dataOut[1916]),
.io_parallelOut_1917(dataOut[1917]),
.io_parallelOut_1918(dataOut[1918]),
.io_parallelOut_1919(dataOut[1919]),
.io_parallelOut_1920(dataOut[1920]),
.io_parallelOut_1921(dataOut[1921]),
.io_parallelOut_1922(dataOut[1922]),
.io_parallelOut_1923(dataOut[1923]),
.io_parallelOut_1924(dataOut[1924]),
.io_parallelOut_1925(dataOut[1925]),
.io_parallelOut_1926(dataOut[1926]),
.io_parallelOut_1927(dataOut[1927]),
.io_parallelOut_1928(dataOut[1928]),
.io_parallelOut_1929(dataOut[1929]),
.io_parallelOut_1930(dataOut[1930]),
.io_parallelOut_1931(dataOut[1931]),
.io_parallelOut_1932(dataOut[1932]),
.io_parallelOut_1933(dataOut[1933]),
.io_parallelOut_1934(dataOut[1934]),
.io_parallelOut_1935(dataOut[1935]),
.io_parallelOut_1936(dataOut[1936]),
.io_parallelOut_1937(dataOut[1937]),
.io_parallelOut_1938(dataOut[1938]),
.io_parallelOut_1939(dataOut[1939]),
.io_parallelOut_1940(dataOut[1940]),
.io_parallelOut_1941(dataOut[1941]),
.io_parallelOut_1942(dataOut[1942]),
.io_parallelOut_1943(dataOut[1943]),
.io_parallelOut_1944(dataOut[1944]),
.io_parallelOut_1945(dataOut[1945]),
.io_parallelOut_1946(dataOut[1946]),
.io_parallelOut_1947(dataOut[1947]),
.io_parallelOut_1948(dataOut[1948]),
.io_parallelOut_1949(dataOut[1949]),
.io_parallelOut_1950(dataOut[1950]),
.io_parallelOut_1951(dataOut[1951]),
.io_parallelOut_1952(dataOut[1952]),
.io_parallelOut_1953(dataOut[1953]),
.io_parallelOut_1954(dataOut[1954]),
.io_parallelOut_1955(dataOut[1955]),
.io_parallelOut_1956(dataOut[1956]),
.io_parallelOut_1957(dataOut[1957]),
.io_parallelOut_1958(dataOut[1958]),
.io_parallelOut_1959(dataOut[1959]),
.io_parallelOut_1960(dataOut[1960]),
.io_parallelOut_1961(dataOut[1961]),
.io_parallelOut_1962(dataOut[1962]),
.io_parallelOut_1963(dataOut[1963]),
.io_parallelOut_1964(dataOut[1964]),
.io_parallelOut_1965(dataOut[1965]),
.io_parallelOut_1966(dataOut[1966]),
.io_parallelOut_1967(dataOut[1967]),
.io_parallelOut_1968(dataOut[1968]),
.io_parallelOut_1969(dataOut[1969]),
.io_parallelOut_1970(dataOut[1970]),
.io_parallelOut_1971(dataOut[1971]),
.io_parallelOut_1972(dataOut[1972]),
.io_parallelOut_1973(dataOut[1973]),
.io_parallelOut_1974(dataOut[1974]),
.io_parallelOut_1975(dataOut[1975]),
.io_parallelOut_1976(dataOut[1976]),
.io_parallelOut_1977(dataOut[1977]),
.io_parallelOut_1978(dataOut[1978]),
.io_parallelOut_1979(dataOut[1979]),
.io_parallelOut_1980(dataOut[1980]),
.io_parallelOut_1981(dataOut[1981]),
.io_parallelOut_1982(dataOut[1982]),
.io_parallelOut_1983(dataOut[1983]),
.io_parallelOut_1984(dataOut[1984]),
.io_parallelOut_1985(dataOut[1985]),
.io_parallelOut_1986(dataOut[1986]),
.io_parallelOut_1987(dataOut[1987]),
.io_parallelOut_1988(dataOut[1988]),
.io_parallelOut_1989(dataOut[1989]),
.io_parallelOut_1990(dataOut[1990]),
.io_parallelOut_1991(dataOut[1991]),
.io_parallelOut_1992(dataOut[1992]),
.io_parallelOut_1993(dataOut[1993]),
.io_parallelOut_1994(dataOut[1994]),
.io_parallelOut_1995(dataOut[1995]),
.io_parallelOut_1996(dataOut[1996]),
.io_parallelOut_1997(dataOut[1997]),
.io_parallelOut_1998(dataOut[1998]),
.io_parallelOut_1999(dataOut[1999]),
.io_parallelOut_2000(dataOut[2000]),
.io_parallelOut_2001(dataOut[2001]),
.io_parallelOut_2002(dataOut[2002]),
.io_parallelOut_2003(dataOut[2003]),
.io_parallelOut_2004(dataOut[2004]),
.io_parallelOut_2005(dataOut[2005]),
.io_parallelOut_2006(dataOut[2006]),
.io_parallelOut_2007(dataOut[2007]),
.io_parallelOut_2008(dataOut[2008]),
.io_parallelOut_2009(dataOut[2009]),
.io_parallelOut_2010(dataOut[2010]),
.io_parallelOut_2011(dataOut[2011]),
.io_parallelOut_2012(dataOut[2012]),
.io_parallelOut_2013(dataOut[2013]),
.io_parallelOut_2014(dataOut[2014]),
.io_parallelOut_2015(dataOut[2015]),
.io_parallelOut_2016(dataOut[2016]),
.io_parallelOut_2017(dataOut[2017]),
.io_parallelOut_2018(dataOut[2018]),
.io_parallelOut_2019(dataOut[2019]),
.io_parallelOut_2020(dataOut[2020]),
.io_parallelOut_2021(dataOut[2021]),
.io_parallelOut_2022(dataOut[2022]),
.io_parallelOut_2023(dataOut[2023]),
.io_parallelOut_2024(dataOut[2024]),
.io_parallelOut_2025(dataOut[2025]),
.io_parallelOut_2026(dataOut[2026]),
.io_parallelOut_2027(dataOut[2027]),
.io_parallelOut_2028(dataOut[2028]),
.io_parallelOut_2029(dataOut[2029]),
.io_parallelOut_2030(dataOut[2030]),
.io_parallelOut_2031(dataOut[2031]),
.io_parallelOut_2032(dataOut[2032]),
.io_parallelOut_2033(dataOut[2033]),
.io_parallelOut_2034(dataOut[2034]),
.io_parallelOut_2035(dataOut[2035]),
.io_parallelOut_2036(dataOut[2036]),
.io_parallelOut_2037(dataOut[2037]),
.io_parallelOut_2038(dataOut[2038]),
.io_parallelOut_2039(dataOut[2039]),
.io_parallelOut_2040(dataOut[2040]),
.io_parallelOut_2041(dataOut[2041]),
.io_parallelOut_2042(dataOut[2042]),
.io_parallelOut_2043(dataOut[2043]),
.io_parallelOut_2044(dataOut[2044]),
.io_parallelOut_2045(dataOut[2045]),
.io_parallelOut_2046(dataOut[2046]),
.io_parallelOut_2047(dataOut[2047]),
.io_parallelOut_2048(dataOut[2048]),
.io_parallelOut_2049(dataOut[2049]),
.io_parallelOut_2050(dataOut[2050]),
.io_parallelOut_2051(dataOut[2051]),
.io_parallelOut_2052(dataOut[2052]),
.io_parallelOut_2053(dataOut[2053]),
.io_parallelOut_2054(dataOut[2054]),
.io_parallelOut_2055(dataOut[2055]),
.io_parallelOut_2056(dataOut[2056]),
.io_parallelOut_2057(dataOut[2057]),
.io_parallelOut_2058(dataOut[2058]),
.io_parallelOut_2059(dataOut[2059]),
.io_parallelOut_2060(dataOut[2060]),
.io_parallelOut_2061(dataOut[2061]),
.io_parallelOut_2062(dataOut[2062]),
.io_parallelOut_2063(dataOut[2063]),
.io_parallelOut_2064(dataOut[2064]),
.io_parallelOut_2065(dataOut[2065]),
.io_parallelOut_2066(dataOut[2066]),
.io_parallelOut_2067(dataOut[2067]),
.io_parallelOut_2068(dataOut[2068]),
.io_parallelOut_2069(dataOut[2069]),
.io_parallelOut_2070(dataOut[2070]),
.io_parallelOut_2071(dataOut[2071]),
.io_parallelOut_2072(dataOut[2072]),
.io_parallelOut_2073(dataOut[2073]),
.io_parallelOut_2074(dataOut[2074]),
.io_parallelOut_2075(dataOut[2075]),
.io_parallelOut_2076(dataOut[2076]),
.io_parallelOut_2077(dataOut[2077]),
.io_parallelOut_2078(dataOut[2078]),
.io_parallelOut_2079(dataOut[2079]),
.io_parallelOut_2080(dataOut[2080]),
.io_parallelOut_2081(dataOut[2081]),
.io_parallelOut_2082(dataOut[2082]),
.io_parallelOut_2083(dataOut[2083]),
.io_parallelOut_2084(dataOut[2084]),
.io_parallelOut_2085(dataOut[2085]),
.io_parallelOut_2086(dataOut[2086]),
.io_parallelOut_2087(dataOut[2087]),
.io_parallelOut_2088(dataOut[2088]),
.io_parallelOut_2089(dataOut[2089]),
.io_parallelOut_2090(dataOut[2090]),
.io_parallelOut_2091(dataOut[2091]),
.io_parallelOut_2092(dataOut[2092]),
.io_parallelOut_2093(dataOut[2093]),
.io_parallelOut_2094(dataOut[2094]),
.io_parallelOut_2095(dataOut[2095]),
.io_parallelOut_2096(dataOut[2096]),
.io_parallelOut_2097(dataOut[2097]),
.io_parallelOut_2098(dataOut[2098]),
.io_parallelOut_2099(dataOut[2099]),
.io_parallelOut_2100(dataOut[2100]),
.io_parallelOut_2101(dataOut[2101]),
.io_parallelOut_2102(dataOut[2102]),
.io_parallelOut_2103(dataOut[2103]),
.io_parallelOut_2104(dataOut[2104]),
.io_parallelOut_2105(dataOut[2105]),
.io_parallelOut_2106(dataOut[2106]),
.io_parallelOut_2107(dataOut[2107]),
.io_parallelOut_2108(dataOut[2108]),
.io_parallelOut_2109(dataOut[2109]),
.io_parallelOut_2110(dataOut[2110]),
.io_parallelOut_2111(dataOut[2111]),
.io_parallelOut_2112(dataOut[2112]),
.io_parallelOut_2113(dataOut[2113]),
.io_parallelOut_2114(dataOut[2114]),
.io_parallelOut_2115(dataOut[2115]),
.io_parallelOut_2116(dataOut[2116]),
.io_parallelOut_2117(dataOut[2117]),
.io_parallelOut_2118(dataOut[2118]),
.io_parallelOut_2119(dataOut[2119]),
.io_parallelOut_2120(dataOut[2120]),
.io_parallelOut_2121(dataOut[2121]),
.io_parallelOut_2122(dataOut[2122]),
.io_parallelOut_2123(dataOut[2123]),
.io_parallelOut_2124(dataOut[2124]),
.io_parallelOut_2125(dataOut[2125]),
.io_parallelOut_2126(dataOut[2126]),
.io_parallelOut_2127(dataOut[2127]),
.io_parallelOut_2128(dataOut[2128]),
.io_parallelOut_2129(dataOut[2129]),
.io_parallelOut_2130(dataOut[2130]),
.io_parallelOut_2131(dataOut[2131]),
.io_parallelOut_2132(dataOut[2132]),
.io_parallelOut_2133(dataOut[2133]),
.io_parallelOut_2134(dataOut[2134]),
.io_parallelOut_2135(dataOut[2135]),
.io_parallelOut_2136(dataOut[2136]),
.io_parallelOut_2137(dataOut[2137]),
.io_parallelOut_2138(dataOut[2138]),
.io_parallelOut_2139(dataOut[2139]),
.io_parallelOut_2140(dataOut[2140]),
.io_parallelOut_2141(dataOut[2141]),
.io_parallelOut_2142(dataOut[2142]),
.io_parallelOut_2143(dataOut[2143]),
.io_parallelOut_2144(dataOut[2144]),
.io_parallelOut_2145(dataOut[2145]),
.io_parallelOut_2146(dataOut[2146]),
.io_parallelOut_2147(dataOut[2147]),
.io_parallelOut_2148(dataOut[2148]),
.io_parallelOut_2149(dataOut[2149]),
.io_parallelOut_2150(dataOut[2150]),
.io_parallelOut_2151(dataOut[2151]),
.io_parallelOut_2152(dataOut[2152]),
.io_parallelOut_2153(dataOut[2153]),
.io_parallelOut_2154(dataOut[2154]),
.io_parallelOut_2155(dataOut[2155]),
.io_parallelOut_2156(dataOut[2156]),
.io_parallelOut_2157(dataOut[2157]),
.io_parallelOut_2158(dataOut[2158]),
.io_parallelOut_2159(dataOut[2159]),
.io_parallelOut_2160(dataOut[2160]),
.io_parallelOut_2161(dataOut[2161]),
.io_parallelOut_2162(dataOut[2162]),
.io_parallelOut_2163(dataOut[2163]),
.io_parallelOut_2164(dataOut[2164]),
.io_parallelOut_2165(dataOut[2165]),
.io_parallelOut_2166(dataOut[2166]),
.io_parallelOut_2167(dataOut[2167]),
.io_parallelOut_2168(dataOut[2168]),
.io_parallelOut_2169(dataOut[2169]),
.io_parallelOut_2170(dataOut[2170]),
.io_parallelOut_2171(dataOut[2171]),
.io_parallelOut_2172(dataOut[2172]),
.io_parallelOut_2173(dataOut[2173]),
.io_parallelOut_2174(dataOut[2174]),
.io_parallelOut_2175(dataOut[2175]),
.io_parallelOut_2176(dataOut[2176]),
.io_parallelOut_2177(dataOut[2177]),
.io_parallelOut_2178(dataOut[2178]),
.io_parallelOut_2179(dataOut[2179]),
.io_parallelOut_2180(dataOut[2180]),
.io_parallelOut_2181(dataOut[2181]),
.io_parallelOut_2182(dataOut[2182]),
.io_parallelOut_2183(dataOut[2183]),
.io_parallelOut_2184(dataOut[2184]),
.io_parallelOut_2185(dataOut[2185]),
.io_parallelOut_2186(dataOut[2186]),
.io_parallelOut_2187(dataOut[2187]),
.io_parallelOut_2188(dataOut[2188]),
.io_parallelOut_2189(dataOut[2189]),
.io_parallelOut_2190(dataOut[2190]),
.io_parallelOut_2191(dataOut[2191]),
.io_parallelOut_2192(dataOut[2192]),
.io_parallelOut_2193(dataOut[2193]),
.io_parallelOut_2194(dataOut[2194]),
.io_parallelOut_2195(dataOut[2195]),
.io_parallelOut_2196(dataOut[2196]),
.io_parallelOut_2197(dataOut[2197]),
.io_parallelOut_2198(dataOut[2198]),
.io_parallelOut_2199(dataOut[2199]),
.io_parallelOut_2200(dataOut[2200]),
.io_parallelOut_2201(dataOut[2201]),
.io_parallelOut_2202(dataOut[2202]),
.io_parallelOut_2203(dataOut[2203]),
.io_parallelOut_2204(dataOut[2204]),
.io_parallelOut_2205(dataOut[2205]),
.io_parallelOut_2206(dataOut[2206]),
.io_parallelOut_2207(dataOut[2207]),
.io_parallelOut_2208(dataOut[2208]),
.io_parallelOut_2209(dataOut[2209]),
.io_parallelOut_2210(dataOut[2210]),
.io_parallelOut_2211(dataOut[2211]),
.io_parallelOut_2212(dataOut[2212]),
.io_parallelOut_2213(dataOut[2213]),
.io_parallelOut_2214(dataOut[2214]),
.io_parallelOut_2215(dataOut[2215]),
.io_parallelOut_2216(dataOut[2216]),
.io_parallelOut_2217(dataOut[2217]),
.io_parallelOut_2218(dataOut[2218]),
.io_parallelOut_2219(dataOut[2219]),
.io_parallelOut_2220(dataOut[2220]),
.io_parallelOut_2221(dataOut[2221]),
.io_parallelOut_2222(dataOut[2222]),
.io_parallelOut_2223(dataOut[2223]),
.io_parallelOut_2224(dataOut[2224]),
.io_parallelOut_2225(dataOut[2225]),
.io_parallelOut_2226(dataOut[2226]),
.io_parallelOut_2227(dataOut[2227]),
.io_parallelOut_2228(dataOut[2228]),
.io_parallelOut_2229(dataOut[2229]),
.io_parallelOut_2230(dataOut[2230]),
.io_parallelOut_2231(dataOut[2231]),
.io_parallelOut_2232(dataOut[2232]),
.io_parallelOut_2233(dataOut[2233]),
.io_parallelOut_2234(dataOut[2234]),
.io_parallelOut_2235(dataOut[2235]),
.io_parallelOut_2236(dataOut[2236]),
.io_parallelOut_2237(dataOut[2237]),
.io_parallelOut_2238(dataOut[2238]),
.io_parallelOut_2239(dataOut[2239]),
.io_parallelOut_2240(dataOut[2240]),
.io_parallelOut_2241(dataOut[2241]),
.io_parallelOut_2242(dataOut[2242]),
.io_parallelOut_2243(dataOut[2243]),
.io_parallelOut_2244(dataOut[2244]),
.io_parallelOut_2245(dataOut[2245]),
.io_parallelOut_2246(dataOut[2246]),
.io_parallelOut_2247(dataOut[2247]),
.io_parallelOut_2248(dataOut[2248]),
.io_parallelOut_2249(dataOut[2249]),
.io_parallelOut_2250(dataOut[2250]),
.io_parallelOut_2251(dataOut[2251]),
.io_parallelOut_2252(dataOut[2252]),
.io_parallelOut_2253(dataOut[2253]),
.io_parallelOut_2254(dataOut[2254]),
.io_parallelOut_2255(dataOut[2255]),
.io_parallelOut_2256(dataOut[2256]),
.io_parallelOut_2257(dataOut[2257]),
.io_parallelOut_2258(dataOut[2258]),
.io_parallelOut_2259(dataOut[2259]),
.io_parallelOut_2260(dataOut[2260]),
.io_parallelOut_2261(dataOut[2261]),
.io_parallelOut_2262(dataOut[2262]),
.io_parallelOut_2263(dataOut[2263]),
.io_parallelOut_2264(dataOut[2264]),
.io_parallelOut_2265(dataOut[2265]),
.io_parallelOut_2266(dataOut[2266]),
.io_parallelOut_2267(dataOut[2267]),
.io_parallelOut_2268(dataOut[2268]),
.io_parallelOut_2269(dataOut[2269]),
.io_parallelOut_2270(dataOut[2270]),
.io_parallelOut_2271(dataOut[2271]),
.io_parallelOut_2272(dataOut[2272]),
.io_parallelOut_2273(dataOut[2273]),
.io_parallelOut_2274(dataOut[2274]),
.io_parallelOut_2275(dataOut[2275]),
.io_parallelOut_2276(dataOut[2276]),
.io_parallelOut_2277(dataOut[2277]),
.io_parallelOut_2278(dataOut[2278]),
.io_parallelOut_2279(dataOut[2279]),
.io_parallelOut_2280(dataOut[2280]),
.io_parallelOut_2281(dataOut[2281]),
.io_parallelOut_2282(dataOut[2282]),
.io_parallelOut_2283(dataOut[2283]),
.io_parallelOut_2284(dataOut[2284]),
.io_parallelOut_2285(dataOut[2285]),
.io_parallelOut_2286(dataOut[2286]),
.io_parallelOut_2287(dataOut[2287]),
.io_parallelOut_2288(dataOut[2288]),
.io_parallelOut_2289(dataOut[2289]),
.io_parallelOut_2290(dataOut[2290]),
.io_parallelOut_2291(dataOut[2291]),
.io_parallelOut_2292(dataOut[2292]),
.io_parallelOut_2293(dataOut[2293]),
.io_parallelOut_2294(dataOut[2294]),
.io_parallelOut_2295(dataOut[2295]),
.io_parallelOut_2296(dataOut[2296]),
.io_parallelOut_2297(dataOut[2297]),
.io_parallelOut_2298(dataOut[2298]),
.io_parallelOut_2299(dataOut[2299]),
.io_parallelOut_2300(dataOut[2300]),
.io_parallelOut_2301(dataOut[2301]),
.io_parallelOut_2302(dataOut[2302]),
.io_parallelOut_2303(dataOut[2303]),
.io_parallelOut_2304(dataOut[2304]),
.io_parallelOut_2305(dataOut[2305]),
.io_parallelOut_2306(dataOut[2306]),
.io_parallelOut_2307(dataOut[2307]),
.io_parallelOut_2308(dataOut[2308]),
.io_parallelOut_2309(dataOut[2309]),
.io_parallelOut_2310(dataOut[2310]),
.io_parallelOut_2311(dataOut[2311]),
.io_parallelOut_2312(dataOut[2312]),
.io_parallelOut_2313(dataOut[2313]),
.io_parallelOut_2314(dataOut[2314]),
.io_parallelOut_2315(dataOut[2315]),
.io_parallelOut_2316(dataOut[2316]),
.io_parallelOut_2317(dataOut[2317]),
.io_parallelOut_2318(dataOut[2318]),
.io_parallelOut_2319(dataOut[2319]),
.io_parallelOut_2320(dataOut[2320]),
.io_parallelOut_2321(dataOut[2321]),
.io_parallelOut_2322(dataOut[2322]),
.io_parallelOut_2323(dataOut[2323]),
.io_parallelOut_2324(dataOut[2324]),
.io_parallelOut_2325(dataOut[2325]),
.io_parallelOut_2326(dataOut[2326]),
.io_parallelOut_2327(dataOut[2327]),
.io_parallelOut_2328(dataOut[2328]),
.io_parallelOut_2329(dataOut[2329]),
.io_parallelOut_2330(dataOut[2330]),
.io_parallelOut_2331(dataOut[2331]),
.io_parallelOut_2332(dataOut[2332]),
.io_parallelOut_2333(dataOut[2333]),
.io_parallelOut_2334(dataOut[2334]),
.io_parallelOut_2335(dataOut[2335]),
.io_parallelOut_2336(dataOut[2336]),
.io_parallelOut_2337(dataOut[2337]),
.io_parallelOut_2338(dataOut[2338]),
.io_parallelOut_2339(dataOut[2339]),
.io_parallelOut_2340(dataOut[2340]),
.io_parallelOut_2341(dataOut[2341]),
.io_parallelOut_2342(dataOut[2342]),
.io_parallelOut_2343(dataOut[2343]),
.io_parallelOut_2344(dataOut[2344]),
.io_parallelOut_2345(dataOut[2345]),
.io_parallelOut_2346(dataOut[2346]),
.io_parallelOut_2347(dataOut[2347]),
.io_parallelOut_2348(dataOut[2348]),
.io_parallelOut_2349(dataOut[2349]),
.io_parallelOut_2350(dataOut[2350]),
.io_parallelOut_2351(dataOut[2351]),
.io_parallelOut_2352(dataOut[2352]),
.io_parallelOut_2353(dataOut[2353]),
.io_parallelOut_2354(dataOut[2354]),
.io_parallelOut_2355(dataOut[2355]),
.io_parallelOut_2356(dataOut[2356]),
.io_parallelOut_2357(dataOut[2357]),
.io_parallelOut_2358(dataOut[2358]),
.io_parallelOut_2359(dataOut[2359]),
.io_parallelOut_2360(dataOut[2360]),
.io_parallelOut_2361(dataOut[2361]),
.io_parallelOut_2362(dataOut[2362]),
.io_parallelOut_2363(dataOut[2363]),
.io_parallelOut_2364(dataOut[2364]),
.io_parallelOut_2365(dataOut[2365]),
.io_parallelOut_2366(dataOut[2366]),
.io_parallelOut_2367(dataOut[2367]),
.io_parallelOut_2368(dataOut[2368]),
.io_parallelOut_2369(dataOut[2369]),
.io_parallelOut_2370(dataOut[2370]),
.io_parallelOut_2371(dataOut[2371]),
.io_parallelOut_2372(dataOut[2372]),
.io_parallelOut_2373(dataOut[2373]),
.io_parallelOut_2374(dataOut[2374]),
.io_parallelOut_2375(dataOut[2375]),
.io_parallelOut_2376(dataOut[2376]),
.io_parallelOut_2377(dataOut[2377]),
.io_parallelOut_2378(dataOut[2378]),
.io_parallelOut_2379(dataOut[2379]),
.io_parallelOut_2380(dataOut[2380]),
.io_parallelOut_2381(dataOut[2381]),
.io_parallelOut_2382(dataOut[2382]),
.io_parallelOut_2383(dataOut[2383]),
.io_parallelOut_2384(dataOut[2384]),
.io_parallelOut_2385(dataOut[2385]),
.io_parallelOut_2386(dataOut[2386]),
.io_parallelOut_2387(dataOut[2387]),
.io_parallelOut_2388(dataOut[2388]),
.io_parallelOut_2389(dataOut[2389]),
.io_parallelOut_2390(dataOut[2390]),
.io_parallelOut_2391(dataOut[2391]),
.io_parallelOut_2392(dataOut[2392]),
.io_parallelOut_2393(dataOut[2393]),
.io_parallelOut_2394(dataOut[2394]),
.io_parallelOut_2395(dataOut[2395]),
.io_parallelOut_2396(dataOut[2396]),
.io_parallelOut_2397(dataOut[2397]),
.io_parallelOut_2398(dataOut[2398]),
.io_parallelOut_2399(dataOut[2399]),
.io_parallelOut_2400(dataOut[2400]),
.io_parallelOut_2401(dataOut[2401]),
.io_parallelOut_2402(dataOut[2402]),
.io_parallelOut_2403(dataOut[2403]),
.io_parallelOut_2404(dataOut[2404]),
.io_parallelOut_2405(dataOut[2405]),
.io_parallelOut_2406(dataOut[2406]),
.io_parallelOut_2407(dataOut[2407]),
.io_parallelOut_2408(dataOut[2408]),
.io_parallelOut_2409(dataOut[2409]),
.io_parallelOut_2410(dataOut[2410]),
.io_parallelOut_2411(dataOut[2411]),
.io_parallelOut_2412(dataOut[2412]),
.io_parallelOut_2413(dataOut[2413]),
.io_parallelOut_2414(dataOut[2414]),
.io_parallelOut_2415(dataOut[2415]),
.io_parallelOut_2416(dataOut[2416]),
.io_parallelOut_2417(dataOut[2417]),
.io_parallelOut_2418(dataOut[2418]),
.io_parallelOut_2419(dataOut[2419]),
.io_parallelOut_2420(dataOut[2420]),
.io_parallelOut_2421(dataOut[2421]),
.io_parallelOut_2422(dataOut[2422]),
.io_parallelOut_2423(dataOut[2423]),
.io_parallelOut_2424(dataOut[2424]),
.io_parallelOut_2425(dataOut[2425]),
.io_parallelOut_2426(dataOut[2426]),
.io_parallelOut_2427(dataOut[2427]),
.io_parallelOut_2428(dataOut[2428]),
.io_parallelOut_2429(dataOut[2429]),
.io_parallelOut_2430(dataOut[2430]),
.io_parallelOut_2431(dataOut[2431]),
.io_parallelOut_2432(dataOut[2432]),
.io_parallelOut_2433(dataOut[2433]),
.io_parallelOut_2434(dataOut[2434]),
.io_parallelOut_2435(dataOut[2435]),
.io_parallelOut_2436(dataOut[2436]),
.io_parallelOut_2437(dataOut[2437]),
.io_parallelOut_2438(dataOut[2438]),
.io_parallelOut_2439(dataOut[2439]),
.io_parallelOut_2440(dataOut[2440]),
.io_parallelOut_2441(dataOut[2441]),
.io_parallelOut_2442(dataOut[2442]),
.io_parallelOut_2443(dataOut[2443]),
.io_parallelOut_2444(dataOut[2444]),
.io_parallelOut_2445(dataOut[2445]),
.io_parallelOut_2446(dataOut[2446]),
.io_parallelOut_2447(dataOut[2447]),
.io_parallelOut_2448(dataOut[2448]),
.io_parallelOut_2449(dataOut[2449]),
.io_parallelOut_2450(dataOut[2450]),
.io_parallelOut_2451(dataOut[2451]),
.io_parallelOut_2452(dataOut[2452]),
.io_parallelOut_2453(dataOut[2453]),
.io_parallelOut_2454(dataOut[2454]),
.io_parallelOut_2455(dataOut[2455]),
.io_parallelOut_2456(dataOut[2456]),
.io_parallelOut_2457(dataOut[2457]),
.io_parallelOut_2458(dataOut[2458]),
.io_parallelOut_2459(dataOut[2459]),
.io_parallelOut_2460(dataOut[2460]),
.io_parallelOut_2461(dataOut[2461]),
.io_parallelOut_2462(dataOut[2462]),
.io_parallelOut_2463(dataOut[2463]),
.io_parallelOut_2464(dataOut[2464]),
.io_parallelOut_2465(dataOut[2465]),
.io_parallelOut_2466(dataOut[2466]),
.io_parallelOut_2467(dataOut[2467]),
.io_parallelOut_2468(dataOut[2468]),
.io_parallelOut_2469(dataOut[2469]),
.io_parallelOut_2470(dataOut[2470]),
.io_parallelOut_2471(dataOut[2471]),
.io_parallelOut_2472(dataOut[2472]),
.io_parallelOut_2473(dataOut[2473]),
.io_parallelOut_2474(dataOut[2474]),
.io_parallelOut_2475(dataOut[2475]),
.io_parallelOut_2476(dataOut[2476]),
.io_parallelOut_2477(dataOut[2477]),
.io_parallelOut_2478(dataOut[2478]),
.io_parallelOut_2479(dataOut[2479]),
.io_parallelOut_2480(dataOut[2480]),
.io_parallelOut_2481(dataOut[2481]),
.io_parallelOut_2482(dataOut[2482]),
.io_parallelOut_2483(dataOut[2483]),
.io_parallelOut_2484(dataOut[2484]),
.io_parallelOut_2485(dataOut[2485]),
.io_parallelOut_2486(dataOut[2486]),
.io_parallelOut_2487(dataOut[2487]),
.io_parallelOut_2488(dataOut[2488]),
.io_parallelOut_2489(dataOut[2489]),
.io_parallelOut_2490(dataOut[2490]),
.io_parallelOut_2491(dataOut[2491]),
.io_parallelOut_2492(dataOut[2492]),
.io_parallelOut_2493(dataOut[2493]),
.io_parallelOut_2494(dataOut[2494]),
.io_parallelOut_2495(dataOut[2495]),
.io_parallelOut_2496(dataOut[2496]),
.io_parallelOut_2497(dataOut[2497]),
.io_parallelOut_2498(dataOut[2498]),
.io_parallelOut_2499(dataOut[2499]),
.io_parallelOut_2500(dataOut[2500]),
.io_parallelOut_2501(dataOut[2501]),
.io_parallelOut_2502(dataOut[2502]),
.io_parallelOut_2503(dataOut[2503]),
.io_parallelOut_2504(dataOut[2504]),
.io_parallelOut_2505(dataOut[2505]),
.io_parallelOut_2506(dataOut[2506]),
.io_parallelOut_2507(dataOut[2507]),
.io_parallelOut_2508(dataOut[2508]),
.io_parallelOut_2509(dataOut[2509]),
.io_parallelOut_2510(dataOut[2510]),
.io_parallelOut_2511(dataOut[2511]),
.io_parallelOut_2512(dataOut[2512]),
.io_parallelOut_2513(dataOut[2513]),
.io_parallelOut_2514(dataOut[2514]),
.io_parallelOut_2515(dataOut[2515]),
.io_parallelOut_2516(dataOut[2516]),
.io_parallelOut_2517(dataOut[2517]),
.io_parallelOut_2518(dataOut[2518]),
.io_parallelOut_2519(dataOut[2519]),
.io_parallelOut_2520(dataOut[2520]),
.io_parallelOut_2521(dataOut[2521]),
.io_parallelOut_2522(dataOut[2522]),
.io_parallelOut_2523(dataOut[2523]),
.io_parallelOut_2524(dataOut[2524]),
.io_parallelOut_2525(dataOut[2525]),
.io_parallelOut_2526(dataOut[2526]),
.io_parallelOut_2527(dataOut[2527]),
.io_parallelOut_2528(dataOut[2528]),
.io_parallelOut_2529(dataOut[2529]),
.io_parallelOut_2530(dataOut[2530]),
.io_parallelOut_2531(dataOut[2531]),
.io_parallelOut_2532(dataOut[2532]),
.io_parallelOut_2533(dataOut[2533]),
.io_parallelOut_2534(dataOut[2534]),
.io_parallelOut_2535(dataOut[2535]),
.io_parallelOut_2536(dataOut[2536]),
.io_parallelOut_2537(dataOut[2537]),
.io_parallelOut_2538(dataOut[2538]),
.io_parallelOut_2539(dataOut[2539]),
.io_parallelOut_2540(dataOut[2540]),
.io_parallelOut_2541(dataOut[2541]),
.io_parallelOut_2542(dataOut[2542]),
.io_parallelOut_2543(dataOut[2543]),
.io_parallelOut_2544(dataOut[2544]),
.io_parallelOut_2545(dataOut[2545]),
.io_parallelOut_2546(dataOut[2546]),
.io_parallelOut_2547(dataOut[2547]),
.io_parallelOut_2548(dataOut[2548]),
.io_parallelOut_2549(dataOut[2549]),
.io_parallelOut_2550(dataOut[2550]),
.io_parallelOut_2551(dataOut[2551]),
.io_parallelOut_2552(dataOut[2552]),
.io_parallelOut_2553(dataOut[2553]),
.io_parallelOut_2554(dataOut[2554]),
.io_parallelOut_2555(dataOut[2555]),
.io_parallelOut_2556(dataOut[2556]),
.io_parallelOut_2557(dataOut[2557]),
.io_parallelOut_2558(dataOut[2558]),
.io_parallelOut_2559(dataOut[2559]),
.io_parallelOut_2560(dataOut[2560]),
.io_parallelOut_2561(dataOut[2561]),
.io_parallelOut_2562(dataOut[2562]),
.io_parallelOut_2563(dataOut[2563]),
.io_parallelOut_2564(dataOut[2564]),
.io_parallelOut_2565(dataOut[2565]),
.io_parallelOut_2566(dataOut[2566]),
.io_parallelOut_2567(dataOut[2567]),
.io_parallelOut_2568(dataOut[2568]),
.io_parallelOut_2569(dataOut[2569]),
.io_parallelOut_2570(dataOut[2570]),
.io_parallelOut_2571(dataOut[2571]),
.io_parallelOut_2572(dataOut[2572]),
.io_parallelOut_2573(dataOut[2573]),
.io_parallelOut_2574(dataOut[2574]),
.io_parallelOut_2575(dataOut[2575]),
.io_parallelOut_2576(dataOut[2576]),
.io_parallelOut_2577(dataOut[2577]),
.io_parallelOut_2578(dataOut[2578]),
.io_parallelOut_2579(dataOut[2579]),
.io_parallelOut_2580(dataOut[2580]),
.io_parallelOut_2581(dataOut[2581]),
.io_parallelOut_2582(dataOut[2582]),
.io_parallelOut_2583(dataOut[2583]),
.io_parallelOut_2584(dataOut[2584]),
.io_parallelOut_2585(dataOut[2585]),
.io_parallelOut_2586(dataOut[2586]),
.io_parallelOut_2587(dataOut[2587]),
.io_parallelOut_2588(dataOut[2588]),
.io_parallelOut_2589(dataOut[2589]),
.io_parallelOut_2590(dataOut[2590]),
.io_parallelOut_2591(dataOut[2591]),
.io_parallelOut_2592(dataOut[2592]),
.io_parallelOut_2593(dataOut[2593]),
.io_parallelOut_2594(dataOut[2594]),
.io_parallelOut_2595(dataOut[2595]),
.io_parallelOut_2596(dataOut[2596]),
.io_parallelOut_2597(dataOut[2597]),
.io_parallelOut_2598(dataOut[2598]),
.io_parallelOut_2599(dataOut[2599]),
.io_parallelOut_2600(dataOut[2600]),
.io_parallelOut_2601(dataOut[2601]),
.io_parallelOut_2602(dataOut[2602]),
.io_parallelOut_2603(dataOut[2603]),
.io_parallelOut_2604(dataOut[2604]),
.io_parallelOut_2605(dataOut[2605]),
.io_parallelOut_2606(dataOut[2606]),
.io_parallelOut_2607(dataOut[2607]),
.io_parallelOut_2608(dataOut[2608]),
.io_parallelOut_2609(dataOut[2609]),
.io_parallelOut_2610(dataOut[2610]),
.io_parallelOut_2611(dataOut[2611]),
.io_parallelOut_2612(dataOut[2612]),
.io_parallelOut_2613(dataOut[2613]),
.io_parallelOut_2614(dataOut[2614]),
.io_parallelOut_2615(dataOut[2615]),
.io_parallelOut_2616(dataOut[2616]),
.io_parallelOut_2617(dataOut[2617]),
.io_parallelOut_2618(dataOut[2618]),
.io_parallelOut_2619(dataOut[2619]),
.io_parallelOut_2620(dataOut[2620]),
.io_parallelOut_2621(dataOut[2621]),
.io_parallelOut_2622(dataOut[2622]),
.io_parallelOut_2623(dataOut[2623]),
.io_parallelOut_2624(dataOut[2624]),
.io_parallelOut_2625(dataOut[2625]),
.io_parallelOut_2626(dataOut[2626]),
.io_parallelOut_2627(dataOut[2627]),
.io_parallelOut_2628(dataOut[2628]),
.io_parallelOut_2629(dataOut[2629]),
.io_parallelOut_2630(dataOut[2630]),
.io_parallelOut_2631(dataOut[2631]),
.io_parallelOut_2632(dataOut[2632]),
.io_parallelOut_2633(dataOut[2633]),
.io_parallelOut_2634(dataOut[2634]),
.io_parallelOut_2635(dataOut[2635]),
.io_parallelOut_2636(dataOut[2636]),
.io_parallelOut_2637(dataOut[2637]),
.io_parallelOut_2638(dataOut[2638]),
.io_parallelOut_2639(dataOut[2639]),
.io_parallelOut_2640(dataOut[2640]),
.io_parallelOut_2641(dataOut[2641]),
.io_parallelOut_2642(dataOut[2642]),
.io_parallelOut_2643(dataOut[2643]),
.io_parallelOut_2644(dataOut[2644]),
.io_parallelOut_2645(dataOut[2645]),
.io_parallelOut_2646(dataOut[2646]),
.io_parallelOut_2647(dataOut[2647]),
.io_parallelOut_2648(dataOut[2648]),
.io_parallelOut_2649(dataOut[2649]),
.io_parallelOut_2650(dataOut[2650]),
.io_parallelOut_2651(dataOut[2651]),
.io_parallelOut_2652(dataOut[2652]),
.io_parallelOut_2653(dataOut[2653]),
.io_parallelOut_2654(dataOut[2654]),
.io_parallelOut_2655(dataOut[2655]),
.io_parallelOut_2656(dataOut[2656]),
.io_parallelOut_2657(dataOut[2657]),
.io_parallelOut_2658(dataOut[2658]),
.io_parallelOut_2659(dataOut[2659]),
.io_parallelOut_2660(dataOut[2660]),
.io_parallelOut_2661(dataOut[2661]),
.io_parallelOut_2662(dataOut[2662]),
.io_parallelOut_2663(dataOut[2663]),
.io_parallelOut_2664(dataOut[2664]),
.io_parallelOut_2665(dataOut[2665]),
.io_parallelOut_2666(dataOut[2666]),
.io_parallelOut_2667(dataOut[2667]),
.io_parallelOut_2668(dataOut[2668]),
.io_parallelOut_2669(dataOut[2669]),
.io_parallelOut_2670(dataOut[2670]),
.io_parallelOut_2671(dataOut[2671]),
.io_parallelOut_2672(dataOut[2672]),
.io_parallelOut_2673(dataOut[2673]),
.io_parallelOut_2674(dataOut[2674]),
.io_parallelOut_2675(dataOut[2675]),
.io_parallelOut_2676(dataOut[2676]),
.io_parallelOut_2677(dataOut[2677]),
.io_parallelOut_2678(dataOut[2678]),
.io_parallelOut_2679(dataOut[2679]),
.io_parallelOut_2680(dataOut[2680]),
.io_parallelOut_2681(dataOut[2681]),
.io_parallelOut_2682(dataOut[2682]),
.io_parallelOut_2683(dataOut[2683]),
.io_parallelOut_2684(dataOut[2684]),
.io_parallelOut_2685(dataOut[2685]),
.io_parallelOut_2686(dataOut[2686]),
.io_parallelOut_2687(dataOut[2687]),
.io_parallelOut_2688(dataOut[2688]),
.io_parallelOut_2689(dataOut[2689]),
.io_parallelOut_2690(dataOut[2690]),
.io_parallelOut_2691(dataOut[2691]),
.io_parallelOut_2692(dataOut[2692]),
.io_parallelOut_2693(dataOut[2693]),
.io_parallelOut_2694(dataOut[2694]),
.io_parallelOut_2695(dataOut[2695]),
.io_parallelOut_2696(dataOut[2696]),
.io_parallelOut_2697(dataOut[2697]),
.io_parallelOut_2698(dataOut[2698]),
.io_parallelOut_2699(dataOut[2699]),
.io_parallelOut_2700(dataOut[2700]),
.io_parallelOut_2701(dataOut[2701]),
.io_parallelOut_2702(dataOut[2702]),
.io_parallelOut_2703(dataOut[2703]),
.io_parallelOut_2704(dataOut[2704]),
.io_parallelOut_2705(dataOut[2705]),
.io_parallelOut_2706(dataOut[2706]),
.io_parallelOut_2707(dataOut[2707]),
.io_parallelOut_2708(dataOut[2708]),
.io_parallelOut_2709(dataOut[2709]),
.io_parallelOut_2710(dataOut[2710]),
.io_parallelOut_2711(dataOut[2711]),
.io_parallelOut_2712(dataOut[2712]),
.io_parallelOut_2713(dataOut[2713]),
.io_parallelOut_2714(dataOut[2714]),
.io_parallelOut_2715(dataOut[2715]),
.io_parallelOut_2716(dataOut[2716]),
.io_parallelOut_2717(dataOut[2717]),
.io_parallelOut_2718(dataOut[2718]),
.io_parallelOut_2719(dataOut[2719]),
.io_parallelOut_2720(dataOut[2720]),
.io_parallelOut_2721(dataOut[2721]),
.io_parallelOut_2722(dataOut[2722]),
.io_parallelOut_2723(dataOut[2723]),
.io_parallelOut_2724(dataOut[2724]),
.io_parallelOut_2725(dataOut[2725]),
.io_parallelOut_2726(dataOut[2726]),
.io_parallelOut_2727(dataOut[2727]),
.io_parallelOut_2728(dataOut[2728]),
.io_parallelOut_2729(dataOut[2729]),
.io_parallelOut_2730(dataOut[2730]),
.io_parallelOut_2731(dataOut[2731]),
.io_parallelOut_2732(dataOut[2732]),
.io_parallelOut_2733(dataOut[2733]),
.io_parallelOut_2734(dataOut[2734]),
.io_parallelOut_2735(dataOut[2735]),
.io_parallelOut_2736(dataOut[2736]),
.io_parallelOut_2737(dataOut[2737]),
.io_parallelOut_2738(dataOut[2738]),
.io_parallelOut_2739(dataOut[2739]),
.io_parallelOut_2740(dataOut[2740]),
.io_parallelOut_2741(dataOut[2741]),
.io_parallelOut_2742(dataOut[2742]),
.io_parallelOut_2743(dataOut[2743]),
.io_parallelOut_2744(dataOut[2744]),
.io_parallelOut_2745(dataOut[2745]),
.io_parallelOut_2746(dataOut[2746]),
.io_parallelOut_2747(dataOut[2747]),
.io_parallelOut_2748(dataOut[2748]),
.io_parallelOut_2749(dataOut[2749]),
.io_parallelOut_2750(dataOut[2750]),
.io_parallelOut_2751(dataOut[2751]),
.io_parallelOut_2752(dataOut[2752]),
.io_parallelOut_2753(dataOut[2753]),
.io_parallelOut_2754(dataOut[2754]),
.io_parallelOut_2755(dataOut[2755]),
.io_parallelOut_2756(dataOut[2756]),
.io_parallelOut_2757(dataOut[2757]),
.io_parallelOut_2758(dataOut[2758]),
.io_parallelOut_2759(dataOut[2759]),
.io_parallelOut_2760(dataOut[2760]),
.io_parallelOut_2761(dataOut[2761]),
.io_parallelOut_2762(dataOut[2762]),
.io_parallelOut_2763(dataOut[2763]),
.io_parallelOut_2764(dataOut[2764]),
.io_parallelOut_2765(dataOut[2765]),
.io_parallelOut_2766(dataOut[2766]),
.io_parallelOut_2767(dataOut[2767]),
.io_parallelOut_2768(dataOut[2768]),
.io_parallelOut_2769(dataOut[2769]),
.io_parallelOut_2770(dataOut[2770]),
.io_parallelOut_2771(dataOut[2771]),
.io_parallelOut_2772(dataOut[2772]),
.io_parallelOut_2773(dataOut[2773]),
.io_parallelOut_2774(dataOut[2774]),
.io_parallelOut_2775(dataOut[2775]),
.io_parallelOut_2776(dataOut[2776]),
.io_parallelOut_2777(dataOut[2777]),
.io_parallelOut_2778(dataOut[2778]),
.io_parallelOut_2779(dataOut[2779]),
.io_parallelOut_2780(dataOut[2780]),
.io_parallelOut_2781(dataOut[2781]),
.io_parallelOut_2782(dataOut[2782]),
.io_parallelOut_2783(dataOut[2783]),
.io_parallelOut_2784(dataOut[2784]),
.io_parallelOut_2785(dataOut[2785]),
.io_parallelOut_2786(dataOut[2786]),
.io_parallelOut_2787(dataOut[2787]),
.io_parallelOut_2788(dataOut[2788]),
.io_parallelOut_2789(dataOut[2789]),
.io_parallelOut_2790(dataOut[2790]),
.io_parallelOut_2791(dataOut[2791]),
.io_parallelOut_2792(dataOut[2792]),
.io_parallelOut_2793(dataOut[2793]),
.io_parallelOut_2794(dataOut[2794]),
.io_parallelOut_2795(dataOut[2795]),
.io_parallelOut_2796(dataOut[2796]),
.io_parallelOut_2797(dataOut[2797]),
.io_parallelOut_2798(dataOut[2798]),
.io_parallelOut_2799(dataOut[2799]),
.io_parallelOut_2800(dataOut[2800]),
.io_parallelOut_2801(dataOut[2801]),
.io_parallelOut_2802(dataOut[2802]),
.io_parallelOut_2803(dataOut[2803]),
.io_parallelOut_2804(dataOut[2804]),
.io_parallelOut_2805(dataOut[2805]),
.io_parallelOut_2806(dataOut[2806]),
.io_parallelOut_2807(dataOut[2807]),
.io_parallelOut_2808(dataOut[2808]),
.io_parallelOut_2809(dataOut[2809]),
.io_parallelOut_2810(dataOut[2810]),
.io_parallelOut_2811(dataOut[2811]),
.io_parallelOut_2812(dataOut[2812]),
.io_parallelOut_2813(dataOut[2813]),
.io_parallelOut_2814(dataOut[2814]),
.io_parallelOut_2815(dataOut[2815]),
.io_parallelOut_2816(dataOut[2816]),
.io_parallelOut_2817(dataOut[2817]),
.io_parallelOut_2818(dataOut[2818]),
.io_parallelOut_2819(dataOut[2819]),
.io_parallelOut_2820(dataOut[2820]),
.io_parallelOut_2821(dataOut[2821]),
.io_parallelOut_2822(dataOut[2822]),
.io_parallelOut_2823(dataOut[2823]),
.io_parallelOut_2824(dataOut[2824]),
.io_parallelOut_2825(dataOut[2825]),
.io_parallelOut_2826(dataOut[2826]),
.io_parallelOut_2827(dataOut[2827]),
.io_parallelOut_2828(dataOut[2828]),
.io_parallelOut_2829(dataOut[2829]),
.io_parallelOut_2830(dataOut[2830]),
.io_parallelOut_2831(dataOut[2831]),
.io_parallelOut_2832(dataOut[2832]),
.io_parallelOut_2833(dataOut[2833]),
.io_parallelOut_2834(dataOut[2834]),
.io_parallelOut_2835(dataOut[2835]),
.io_parallelOut_2836(dataOut[2836]),
.io_parallelOut_2837(dataOut[2837]),
.io_parallelOut_2838(dataOut[2838]),
.io_parallelOut_2839(dataOut[2839]),
.io_parallelOut_2840(dataOut[2840]),
.io_parallelOut_2841(dataOut[2841]),
.io_parallelOut_2842(dataOut[2842]),
.io_parallelOut_2843(dataOut[2843]),
.io_parallelOut_2844(dataOut[2844]),
.io_parallelOut_2845(dataOut[2845]),
.io_parallelOut_2846(dataOut[2846]),
.io_parallelOut_2847(dataOut[2847]),
.io_parallelOut_2848(dataOut[2848]),
.io_parallelOut_2849(dataOut[2849]),
.io_parallelOut_2850(dataOut[2850]),
.io_parallelOut_2851(dataOut[2851]),
.io_parallelOut_2852(dataOut[2852]),
.io_parallelOut_2853(dataOut[2853]),
.io_parallelOut_2854(dataOut[2854]),
.io_parallelOut_2855(dataOut[2855]),
.io_parallelOut_2856(dataOut[2856]),
.io_parallelOut_2857(dataOut[2857]),
.io_parallelOut_2858(dataOut[2858]),
.io_parallelOut_2859(dataOut[2859]),
.io_parallelOut_2860(dataOut[2860]),
.io_parallelOut_2861(dataOut[2861]),
.io_parallelOut_2862(dataOut[2862]),
.io_parallelOut_2863(dataOut[2863]),
.io_parallelOut_2864(dataOut[2864]),
.io_parallelOut_2865(dataOut[2865]),
.io_parallelOut_2866(dataOut[2866]),
.io_parallelOut_2867(dataOut[2867]),
.io_parallelOut_2868(dataOut[2868]),
.io_parallelOut_2869(dataOut[2869]),
.io_parallelOut_2870(dataOut[2870]),
.io_parallelOut_2871(dataOut[2871]),
.io_parallelOut_2872(dataOut[2872]),
.io_parallelOut_2873(dataOut[2873]),
.io_parallelOut_2874(dataOut[2874]),
.io_parallelOut_2875(dataOut[2875]),
.io_parallelOut_2876(dataOut[2876]),
.io_parallelOut_2877(dataOut[2877]),
.io_parallelOut_2878(dataOut[2878]),
.io_parallelOut_2879(dataOut[2879]),
.io_parallelOut_2880(dataOut[2880]),
.io_parallelOut_2881(dataOut[2881]),
.io_parallelOut_2882(dataOut[2882]),
.io_parallelOut_2883(dataOut[2883]),
.io_parallelOut_2884(dataOut[2884]),
.io_parallelOut_2885(dataOut[2885]),
.io_parallelOut_2886(dataOut[2886]),
.io_parallelOut_2887(dataOut[2887]),
.io_parallelOut_2888(dataOut[2888]),
.io_parallelOut_2889(dataOut[2889]),
.io_parallelOut_2890(dataOut[2890]),
.io_parallelOut_2891(dataOut[2891]),
.io_parallelOut_2892(dataOut[2892]),
.io_parallelOut_2893(dataOut[2893]),
.io_parallelOut_2894(dataOut[2894]),
.io_parallelOut_2895(dataOut[2895]),
.io_parallelOut_2896(dataOut[2896]),
.io_parallelOut_2897(dataOut[2897]),
.io_parallelOut_2898(dataOut[2898]),
.io_parallelOut_2899(dataOut[2899]),
.io_parallelOut_2900(dataOut[2900]),
.io_parallelOut_2901(dataOut[2901]),
.io_parallelOut_2902(dataOut[2902]),
.io_parallelOut_2903(dataOut[2903]),
.io_parallelOut_2904(dataOut[2904]),
.io_parallelOut_2905(dataOut[2905]),
.io_parallelOut_2906(dataOut[2906]),
.io_parallelOut_2907(dataOut[2907]),
.io_parallelOut_2908(dataOut[2908]),
.io_parallelOut_2909(dataOut[2909]),
.io_parallelOut_2910(dataOut[2910]),
.io_parallelOut_2911(dataOut[2911]),
.io_parallelOut_2912(dataOut[2912]),
.io_parallelOut_2913(dataOut[2913]),
.io_parallelOut_2914(dataOut[2914]),
.io_parallelOut_2915(dataOut[2915]),
.io_parallelOut_2916(dataOut[2916]),
.io_parallelOut_2917(dataOut[2917]),
.io_parallelOut_2918(dataOut[2918]),
.io_parallelOut_2919(dataOut[2919]),
.io_parallelOut_2920(dataOut[2920]),
.io_parallelOut_2921(dataOut[2921]),
.io_parallelOut_2922(dataOut[2922]),
.io_parallelOut_2923(dataOut[2923]),
.io_parallelOut_2924(dataOut[2924]),
.io_parallelOut_2925(dataOut[2925]),
.io_parallelOut_2926(dataOut[2926]),
.io_parallelOut_2927(dataOut[2927]),
.io_parallelOut_2928(dataOut[2928]),
.io_parallelOut_2929(dataOut[2929]),
.io_parallelOut_2930(dataOut[2930]),
.io_parallelOut_2931(dataOut[2931]),
.io_parallelOut_2932(dataOut[2932]),
.io_parallelOut_2933(dataOut[2933]),
.io_parallelOut_2934(dataOut[2934]),
.io_parallelOut_2935(dataOut[2935]),
.io_parallelOut_2936(dataOut[2936]),
.io_parallelOut_2937(dataOut[2937]),
.io_parallelOut_2938(dataOut[2938]),
.io_parallelOut_2939(dataOut[2939]),
.io_parallelOut_2940(dataOut[2940]),
.io_parallelOut_2941(dataOut[2941]),
.io_parallelOut_2942(dataOut[2942]),
.io_parallelOut_2943(dataOut[2943]),
.io_parallelOut_2944(dataOut[2944]),
.io_parallelOut_2945(dataOut[2945]),
.io_parallelOut_2946(dataOut[2946]),
.io_parallelOut_2947(dataOut[2947]),
.io_parallelOut_2948(dataOut[2948]),
.io_parallelOut_2949(dataOut[2949]),
.io_parallelOut_2950(dataOut[2950]),
.io_parallelOut_2951(dataOut[2951]),
.io_parallelOut_2952(dataOut[2952]),
.io_parallelOut_2953(dataOut[2953]),
.io_parallelOut_2954(dataOut[2954]),
.io_parallelOut_2955(dataOut[2955]),
.io_parallelOut_2956(dataOut[2956]),
.io_parallelOut_2957(dataOut[2957]),
.io_parallelOut_2958(dataOut[2958]),
.io_parallelOut_2959(dataOut[2959]),
.io_parallelOut_2960(dataOut[2960]),
.io_parallelOut_2961(dataOut[2961]),
.io_parallelOut_2962(dataOut[2962]),
.io_parallelOut_2963(dataOut[2963]),
.io_parallelOut_2964(dataOut[2964]),
.io_parallelOut_2965(dataOut[2965]),
.io_parallelOut_2966(dataOut[2966]),
.io_parallelOut_2967(dataOut[2967]),
.io_parallelOut_2968(dataOut[2968]),
.io_parallelOut_2969(dataOut[2969]),
.io_parallelOut_2970(dataOut[2970]),
.io_parallelOut_2971(dataOut[2971]),
.io_parallelOut_2972(dataOut[2972]),
.io_parallelOut_2973(dataOut[2973]),
.io_parallelOut_2974(dataOut[2974]),
.io_parallelOut_2975(dataOut[2975]),
.io_parallelOut_2976(dataOut[2976]),
.io_parallelOut_2977(dataOut[2977]),
.io_parallelOut_2978(dataOut[2978]),
.io_parallelOut_2979(dataOut[2979]),
.io_parallelOut_2980(dataOut[2980]),
.io_parallelOut_2981(dataOut[2981]),
.io_parallelOut_2982(dataOut[2982]),
.io_parallelOut_2983(dataOut[2983]),
.io_parallelOut_2984(dataOut[2984]),
.io_parallelOut_2985(dataOut[2985]),
.io_parallelOut_2986(dataOut[2986]),
.io_parallelOut_2987(dataOut[2987]),
.io_parallelOut_2988(dataOut[2988]),
.io_parallelOut_2989(dataOut[2989]),
.io_parallelOut_2990(dataOut[2990]),
.io_parallelOut_2991(dataOut[2991]),
.io_parallelOut_2992(dataOut[2992]),
.io_parallelOut_2993(dataOut[2993]),
.io_parallelOut_2994(dataOut[2994]),
.io_parallelOut_2995(dataOut[2995]),
.io_parallelOut_2996(dataOut[2996]),
.io_parallelOut_2997(dataOut[2997]),
.io_parallelOut_2998(dataOut[2998]),
.io_parallelOut_2999(dataOut[2999]),
.io_parallelOut_3000(dataOut[3000]),
.io_parallelOut_3001(dataOut[3001]),
.io_parallelOut_3002(dataOut[3002]),
.io_parallelOut_3003(dataOut[3003]),
.io_parallelOut_3004(dataOut[3004]),
.io_parallelOut_3005(dataOut[3005]),
.io_parallelOut_3006(dataOut[3006]),
.io_parallelOut_3007(dataOut[3007]),
.io_parallelOut_3008(dataOut[3008]),
.io_parallelOut_3009(dataOut[3009]),
.io_parallelOut_3010(dataOut[3010]),
.io_parallelOut_3011(dataOut[3011]),
.io_parallelOut_3012(dataOut[3012]),
.io_parallelOut_3013(dataOut[3013]),
.io_parallelOut_3014(dataOut[3014]),
.io_parallelOut_3015(dataOut[3015]),
.io_parallelOut_3016(dataOut[3016]),
.io_parallelOut_3017(dataOut[3017]),
.io_parallelOut_3018(dataOut[3018]),
.io_parallelOut_3019(dataOut[3019]),
.io_parallelOut_3020(dataOut[3020]),
.io_parallelOut_3021(dataOut[3021]),
.io_parallelOut_3022(dataOut[3022]),
.io_parallelOut_3023(dataOut[3023]),
.io_parallelOut_3024(dataOut[3024]),
.io_parallelOut_3025(dataOut[3025]),
.io_parallelOut_3026(dataOut[3026]),
.io_parallelOut_3027(dataOut[3027]),
.io_parallelOut_3028(dataOut[3028]),
.io_parallelOut_3029(dataOut[3029]),
.io_parallelOut_3030(dataOut[3030]),
.io_parallelOut_3031(dataOut[3031]),
.io_parallelOut_3032(dataOut[3032]),
.io_parallelOut_3033(dataOut[3033]),
.io_parallelOut_3034(dataOut[3034]),
.io_parallelOut_3035(dataOut[3035]),
.io_parallelOut_3036(dataOut[3036]),
.io_parallelOut_3037(dataOut[3037]),
.io_parallelOut_3038(dataOut[3038]),
.io_parallelOut_3039(dataOut[3039]),
.io_parallelOut_3040(dataOut[3040]),
.io_parallelOut_3041(dataOut[3041]),
.io_parallelOut_3042(dataOut[3042]),
.io_parallelOut_3043(dataOut[3043]),
.io_parallelOut_3044(dataOut[3044]),
.io_parallelOut_3045(dataOut[3045]),
.io_parallelOut_3046(dataOut[3046]),
.io_parallelOut_3047(dataOut[3047]),
.io_parallelOut_3048(dataOut[3048]),
.io_parallelOut_3049(dataOut[3049]),
.io_parallelOut_3050(dataOut[3050]),
.io_parallelOut_3051(dataOut[3051]),
.io_parallelOut_3052(dataOut[3052]),
.io_parallelOut_3053(dataOut[3053]),
.io_parallelOut_3054(dataOut[3054]),
.io_parallelOut_3055(dataOut[3055]),
.io_parallelOut_3056(dataOut[3056]),
.io_parallelOut_3057(dataOut[3057]),
.io_parallelOut_3058(dataOut[3058]),
.io_parallelOut_3059(dataOut[3059]),
.io_parallelOut_3060(dataOut[3060]),
.io_parallelOut_3061(dataOut[3061]),
.io_parallelOut_3062(dataOut[3062]),
.io_parallelOut_3063(dataOut[3063]),
.io_parallelOut_3064(dataOut[3064]),
.io_parallelOut_3065(dataOut[3065]),
.io_parallelOut_3066(dataOut[3066]),
.io_parallelOut_3067(dataOut[3067]),
.io_parallelOut_3068(dataOut[3068]),
.io_parallelOut_3069(dataOut[3069]),
.io_parallelOut_3070(dataOut[3070]),
.io_parallelOut_3071(dataOut[3071]),
.io_parallelOut_3072(dataOut[3072]),
.io_parallelOut_3073(dataOut[3073]),
.io_parallelOut_3074(dataOut[3074]),
.io_parallelOut_3075(dataOut[3075]),
.io_parallelOut_3076(dataOut[3076]),
.io_parallelOut_3077(dataOut[3077]),
.io_parallelOut_3078(dataOut[3078]),
.io_parallelOut_3079(dataOut[3079]),
.io_parallelOut_3080(dataOut[3080]),
.io_parallelOut_3081(dataOut[3081]),
.io_parallelOut_3082(dataOut[3082]),
.io_parallelOut_3083(dataOut[3083]),
.io_parallelOut_3084(dataOut[3084]),
.io_parallelOut_3085(dataOut[3085]),
.io_parallelOut_3086(dataOut[3086]),
.io_parallelOut_3087(dataOut[3087]),
.io_parallelOut_3088(dataOut[3088]),
.io_parallelOut_3089(dataOut[3089]),
.io_parallelOut_3090(dataOut[3090]),
.io_parallelOut_3091(dataOut[3091]),
.io_parallelOut_3092(dataOut[3092]),
.io_parallelOut_3093(dataOut[3093]),
.io_parallelOut_3094(dataOut[3094]),
.io_parallelOut_3095(dataOut[3095]),
.io_parallelOut_3096(dataOut[3096]),
.io_parallelOut_3097(dataOut[3097]),
.io_parallelOut_3098(dataOut[3098]),
.io_parallelOut_3099(dataOut[3099]),
.io_parallelOut_3100(dataOut[3100]),
.io_parallelOut_3101(dataOut[3101]),
.io_parallelOut_3102(dataOut[3102]),
.io_parallelOut_3103(dataOut[3103]),
.io_parallelOut_3104(dataOut[3104]),
.io_parallelOut_3105(dataOut[3105]),
.io_parallelOut_3106(dataOut[3106]),
.io_parallelOut_3107(dataOut[3107]),
.io_parallelOut_3108(dataOut[3108]),
.io_parallelOut_3109(dataOut[3109]),
.io_parallelOut_3110(dataOut[3110]),
.io_parallelOut_3111(dataOut[3111]),
.io_parallelOut_3112(dataOut[3112]),
.io_parallelOut_3113(dataOut[3113]),
.io_parallelOut_3114(dataOut[3114]),
.io_parallelOut_3115(dataOut[3115]),
.io_parallelOut_3116(dataOut[3116]),
.io_parallelOut_3117(dataOut[3117]),
.io_parallelOut_3118(dataOut[3118]),
.io_parallelOut_3119(dataOut[3119]),
.io_parallelOut_3120(dataOut[3120]),
.io_parallelOut_3121(dataOut[3121]),
.io_parallelOut_3122(dataOut[3122]),
.io_parallelOut_3123(dataOut[3123]),
.io_parallelOut_3124(dataOut[3124]),
.io_parallelOut_3125(dataOut[3125]),
.io_parallelOut_3126(dataOut[3126]),
.io_parallelOut_3127(dataOut[3127]),
.io_parallelOut_3128(dataOut[3128]),
.io_parallelOut_3129(dataOut[3129]),
.io_parallelOut_3130(dataOut[3130]),
.io_parallelOut_3131(dataOut[3131]),
.io_parallelOut_3132(dataOut[3132]),
.io_parallelOut_3133(dataOut[3133]),
.io_parallelOut_3134(dataOut[3134]),
.io_parallelOut_3135(dataOut[3135]),
.io_parallelOut_3136(dataOut[3136]),
.io_parallelOut_3137(dataOut[3137]),
.io_parallelOut_3138(dataOut[3138]),
.io_parallelOut_3139(dataOut[3139]),
.io_parallelOut_3140(dataOut[3140]),
.io_parallelOut_3141(dataOut[3141]),
.io_parallelOut_3142(dataOut[3142]),
.io_parallelOut_3143(dataOut[3143]),
.io_parallelOut_3144(dataOut[3144]),
.io_parallelOut_3145(dataOut[3145]),
.io_parallelOut_3146(dataOut[3146]),
.io_parallelOut_3147(dataOut[3147]),
.io_parallelOut_3148(dataOut[3148]),
.io_parallelOut_3149(dataOut[3149]),
.io_parallelOut_3150(dataOut[3150]),
.io_parallelOut_3151(dataOut[3151]),
.io_parallelOut_3152(dataOut[3152]),
.io_parallelOut_3153(dataOut[3153]),
.io_parallelOut_3154(dataOut[3154]),
.io_parallelOut_3155(dataOut[3155]),
.io_parallelOut_3156(dataOut[3156]),
.io_parallelOut_3157(dataOut[3157]),
.io_parallelOut_3158(dataOut[3158]),
.io_parallelOut_3159(dataOut[3159]),
.io_parallelOut_3160(dataOut[3160]),
.io_parallelOut_3161(dataOut[3161]),
.io_parallelOut_3162(dataOut[3162]),
.io_parallelOut_3163(dataOut[3163]),
.io_parallelOut_3164(dataOut[3164]),
.io_parallelOut_3165(dataOut[3165]),
.io_parallelOut_3166(dataOut[3166]),
.io_parallelOut_3167(dataOut[3167]),
.io_parallelOut_3168(dataOut[3168]),
.io_parallelOut_3169(dataOut[3169]),
.io_parallelOut_3170(dataOut[3170]),
.io_parallelOut_3171(dataOut[3171]),
.io_parallelOut_3172(dataOut[3172]),
.io_parallelOut_3173(dataOut[3173]),
.io_parallelOut_3174(dataOut[3174]),
.io_parallelOut_3175(dataOut[3175]),
.io_parallelOut_3176(dataOut[3176]),
.io_parallelOut_3177(dataOut[3177]),
.io_parallelOut_3178(dataOut[3178]),
.io_parallelOut_3179(dataOut[3179]),
.io_parallelOut_3180(dataOut[3180]),
.io_parallelOut_3181(dataOut[3181]),
.io_parallelOut_3182(dataOut[3182]),
.io_parallelOut_3183(dataOut[3183]),
.io_parallelOut_3184(dataOut[3184]),
.io_parallelOut_3185(dataOut[3185]),
.io_parallelOut_3186(dataOut[3186]),
.io_parallelOut_3187(dataOut[3187]),
.io_parallelOut_3188(dataOut[3188]),
.io_parallelOut_3189(dataOut[3189]),
.io_parallelOut_3190(dataOut[3190]),
.io_parallelOut_3191(dataOut[3191]),
.io_parallelOut_3192(dataOut[3192]),
.io_parallelOut_3193(dataOut[3193]),
.io_parallelOut_3194(dataOut[3194]),
.io_parallelOut_3195(dataOut[3195]),
.io_parallelOut_3196(dataOut[3196]),
.io_parallelOut_3197(dataOut[3197]),
.io_parallelOut_3198(dataOut[3198]),
.io_parallelOut_3199(dataOut[3199]),
.io_parallelOut_3200(dataOut[3200]),
.io_parallelOut_3201(dataOut[3201]),
.io_parallelOut_3202(dataOut[3202]),
.io_parallelOut_3203(dataOut[3203]),
.io_parallelOut_3204(dataOut[3204]),
.io_parallelOut_3205(dataOut[3205]),
.io_parallelOut_3206(dataOut[3206]),
.io_parallelOut_3207(dataOut[3207]),
.io_parallelOut_3208(dataOut[3208]),
.io_parallelOut_3209(dataOut[3209]),
.io_parallelOut_3210(dataOut[3210]),
.io_parallelOut_3211(dataOut[3211]),
.io_parallelOut_3212(dataOut[3212]),
.io_parallelOut_3213(dataOut[3213]),
.io_parallelOut_3214(dataOut[3214]),
.io_parallelOut_3215(dataOut[3215]),
.io_parallelOut_3216(dataOut[3216]),
.io_parallelOut_3217(dataOut[3217]),
.io_parallelOut_3218(dataOut[3218]),
.io_parallelOut_3219(dataOut[3219]),
.io_parallelOut_3220(dataOut[3220]),
.io_parallelOut_3221(dataOut[3221]),
.io_parallelOut_3222(dataOut[3222]),
.io_parallelOut_3223(dataOut[3223]),
.io_parallelOut_3224(dataOut[3224]),
.io_parallelOut_3225(dataOut[3225]),
.io_parallelOut_3226(dataOut[3226]),
.io_parallelOut_3227(dataOut[3227]),
.io_parallelOut_3228(dataOut[3228]),
.io_parallelOut_3229(dataOut[3229]),
.io_parallelOut_3230(dataOut[3230]),
.io_parallelOut_3231(dataOut[3231]),
.io_parallelOut_3232(dataOut[3232]),
.io_parallelOut_3233(dataOut[3233]),
.io_parallelOut_3234(dataOut[3234]),
.io_parallelOut_3235(dataOut[3235]),
.io_parallelOut_3236(dataOut[3236]),
.io_parallelOut_3237(dataOut[3237]),
.io_parallelOut_3238(dataOut[3238]),
.io_parallelOut_3239(dataOut[3239]),
.io_parallelOut_3240(dataOut[3240]),
.io_parallelOut_3241(dataOut[3241]),
.io_parallelOut_3242(dataOut[3242]),
.io_parallelOut_3243(dataOut[3243]),
.io_parallelOut_3244(dataOut[3244]),
.io_parallelOut_3245(dataOut[3245]),
.io_parallelOut_3246(dataOut[3246]),
.io_parallelOut_3247(dataOut[3247]),
.io_parallelOut_3248(dataOut[3248]),
.io_parallelOut_3249(dataOut[3249]),
.io_parallelOut_3250(dataOut[3250]),
.io_parallelOut_3251(dataOut[3251]),
.io_parallelOut_3252(dataOut[3252]),
.io_parallelOut_3253(dataOut[3253]),
.io_parallelOut_3254(dataOut[3254]),
.io_parallelOut_3255(dataOut[3255]),
.io_parallelOut_3256(dataOut[3256]),
.io_parallelOut_3257(dataOut[3257]),
.io_parallelOut_3258(dataOut[3258]),
.io_parallelOut_3259(dataOut[3259]),
.io_parallelOut_3260(dataOut[3260]),
.io_parallelOut_3261(dataOut[3261]),
.io_parallelOut_3262(dataOut[3262]),
.io_parallelOut_3263(dataOut[3263]),
.io_parallelOut_3264(dataOut[3264]),
.io_parallelOut_3265(dataOut[3265]),
.io_parallelOut_3266(dataOut[3266]),
.io_parallelOut_3267(dataOut[3267]),
.io_parallelOut_3268(dataOut[3268]),
.io_parallelOut_3269(dataOut[3269]),
.io_parallelOut_3270(dataOut[3270]),
.io_parallelOut_3271(dataOut[3271]),
.io_parallelOut_3272(dataOut[3272]),
.io_parallelOut_3273(dataOut[3273]),
.io_parallelOut_3274(dataOut[3274]),
.io_parallelOut_3275(dataOut[3275]),
.io_parallelOut_3276(dataOut[3276]),
.io_parallelOut_3277(dataOut[3277]),
.io_parallelOut_3278(dataOut[3278]),
.io_parallelOut_3279(dataOut[3279]),
.io_parallelOut_3280(dataOut[3280]),
.io_parallelOut_3281(dataOut[3281]),
.io_parallelOut_3282(dataOut[3282]),
.io_parallelOut_3283(dataOut[3283]),
.io_parallelOut_3284(dataOut[3284]),
.io_parallelOut_3285(dataOut[3285]),
.io_parallelOut_3286(dataOut[3286]),
.io_parallelOut_3287(dataOut[3287]),
.io_parallelOut_3288(dataOut[3288]),
.io_parallelOut_3289(dataOut[3289]),
.io_parallelOut_3290(dataOut[3290]),
.io_parallelOut_3291(dataOut[3291]),
.io_parallelOut_3292(dataOut[3292]),
.io_parallelOut_3293(dataOut[3293]),
.io_parallelOut_3294(dataOut[3294]),
.io_parallelOut_3295(dataOut[3295]),
.io_parallelOut_3296(dataOut[3296]),
.io_parallelOut_3297(dataOut[3297]),
.io_parallelOut_3298(dataOut[3298]),
.io_parallelOut_3299(dataOut[3299]),
.io_parallelOut_3300(dataOut[3300]),
.io_parallelOut_3301(dataOut[3301]),
.io_parallelOut_3302(dataOut[3302]),
.io_parallelOut_3303(dataOut[3303]),
.io_parallelOut_3304(dataOut[3304]),
.io_parallelOut_3305(dataOut[3305]),
.io_parallelOut_3306(dataOut[3306]),
.io_parallelOut_3307(dataOut[3307]),
.io_parallelOut_3308(dataOut[3308]),
.io_parallelOut_3309(dataOut[3309]),
.io_parallelOut_3310(dataOut[3310]),
.io_parallelOut_3311(dataOut[3311]),
.io_parallelOut_3312(dataOut[3312]),
.io_parallelOut_3313(dataOut[3313]),
.io_parallelOut_3314(dataOut[3314]),
.io_parallelOut_3315(dataOut[3315]),
.io_parallelOut_3316(dataOut[3316]),
.io_parallelOut_3317(dataOut[3317]),
.io_parallelOut_3318(dataOut[3318]),
.io_parallelOut_3319(dataOut[3319]),
.io_parallelOut_3320(dataOut[3320]),
.io_parallelOut_3321(dataOut[3321]),
.io_parallelOut_3322(dataOut[3322]),
.io_parallelOut_3323(dataOut[3323]),
.io_parallelOut_3324(dataOut[3324]),
.io_parallelOut_3325(dataOut[3325]),
.io_parallelOut_3326(dataOut[3326]),
.io_parallelOut_3327(dataOut[3327]),
.io_parallelOut_3328(dataOut[3328]),
.io_parallelOut_3329(dataOut[3329]),
.io_parallelOut_3330(dataOut[3330]),
.io_parallelOut_3331(dataOut[3331]),
.io_parallelOut_3332(dataOut[3332]),
.io_parallelOut_3333(dataOut[3333]),
.io_parallelOut_3334(dataOut[3334]),
.io_parallelOut_3335(dataOut[3335]),
.io_parallelOut_3336(dataOut[3336]),
.io_parallelOut_3337(dataOut[3337]),
.io_parallelOut_3338(dataOut[3338]),
.io_parallelOut_3339(dataOut[3339]),
.io_parallelOut_3340(dataOut[3340]),
.io_parallelOut_3341(dataOut[3341]),
.io_parallelOut_3342(dataOut[3342]),
.io_parallelOut_3343(dataOut[3343]),
.io_parallelOut_3344(dataOut[3344]),
.io_parallelOut_3345(dataOut[3345]),
.io_parallelOut_3346(dataOut[3346]),
.io_parallelOut_3347(dataOut[3347]),
.io_parallelOut_3348(dataOut[3348]),
.io_parallelOut_3349(dataOut[3349]),
.io_parallelOut_3350(dataOut[3350]),
.io_parallelOut_3351(dataOut[3351]),
.io_parallelOut_3352(dataOut[3352]),
.io_parallelOut_3353(dataOut[3353]),
.io_parallelOut_3354(dataOut[3354]),
.io_parallelOut_3355(dataOut[3355]),
.io_parallelOut_3356(dataOut[3356]),
.io_parallelOut_3357(dataOut[3357]),
.io_parallelOut_3358(dataOut[3358]),
.io_parallelOut_3359(dataOut[3359]),
.io_parallelOut_3360(dataOut[3360]),
.io_parallelOut_3361(dataOut[3361]),
.io_parallelOut_3362(dataOut[3362]),
.io_parallelOut_3363(dataOut[3363]),
.io_parallelOut_3364(dataOut[3364]),
.io_parallelOut_3365(dataOut[3365]),
.io_parallelOut_3366(dataOut[3366]),
.io_parallelOut_3367(dataOut[3367]),
.io_parallelOut_3368(dataOut[3368]),
.io_parallelOut_3369(dataOut[3369]),
.io_parallelOut_3370(dataOut[3370]),
.io_parallelOut_3371(dataOut[3371]),
.io_parallelOut_3372(dataOut[3372]),
.io_parallelOut_3373(dataOut[3373]),
.io_parallelOut_3374(dataOut[3374]),
.io_parallelOut_3375(dataOut[3375]),
.io_parallelOut_3376(dataOut[3376]),
.io_parallelOut_3377(dataOut[3377]),
.io_parallelOut_3378(dataOut[3378]),
.io_parallelOut_3379(dataOut[3379]),
.io_parallelOut_3380(dataOut[3380]),
.io_parallelOut_3381(dataOut[3381]),
.io_parallelOut_3382(dataOut[3382]),
.io_parallelOut_3383(dataOut[3383]),
.io_parallelOut_3384(dataOut[3384]),
.io_parallelOut_3385(dataOut[3385]),
.io_parallelOut_3386(dataOut[3386]),
.io_parallelOut_3387(dataOut[3387]),
.io_parallelOut_3388(dataOut[3388]),
.io_parallelOut_3389(dataOut[3389]),
.io_parallelOut_3390(dataOut[3390]),
.io_parallelOut_3391(dataOut[3391]),
.io_parallelOut_3392(dataOut[3392]),
.io_parallelOut_3393(dataOut[3393]),
.io_parallelOut_3394(dataOut[3394]),
.io_parallelOut_3395(dataOut[3395]),
.io_parallelOut_3396(dataOut[3396]),
.io_parallelOut_3397(dataOut[3397]),
.io_parallelOut_3398(dataOut[3398]),
.io_parallelOut_3399(dataOut[3399]),
.io_parallelOut_3400(dataOut[3400]),
.io_parallelOut_3401(dataOut[3401]),
.io_parallelOut_3402(dataOut[3402]),
.io_parallelOut_3403(dataOut[3403]),
.io_parallelOut_3404(dataOut[3404]),
.io_parallelOut_3405(dataOut[3405]),
.io_parallelOut_3406(dataOut[3406]),
.io_parallelOut_3407(dataOut[3407]),
.io_parallelOut_3408(dataOut[3408]),
.io_parallelOut_3409(dataOut[3409]),
.io_parallelOut_3410(dataOut[3410]),
.io_parallelOut_3411(dataOut[3411]),
.io_parallelOut_3412(dataOut[3412]),
.io_parallelOut_3413(dataOut[3413]),
.io_parallelOut_3414(dataOut[3414]),
.io_parallelOut_3415(dataOut[3415]),
.io_parallelOut_3416(dataOut[3416]),
.io_parallelOut_3417(dataOut[3417]),
.io_parallelOut_3418(dataOut[3418]),
.io_parallelOut_3419(dataOut[3419]),
.io_parallelOut_3420(dataOut[3420]),
.io_parallelOut_3421(dataOut[3421]),
.io_parallelOut_3422(dataOut[3422]),
.io_parallelOut_3423(dataOut[3423]),
.io_parallelOut_3424(dataOut[3424]),
.io_parallelOut_3425(dataOut[3425]),
.io_parallelOut_3426(dataOut[3426]),
.io_parallelOut_3427(dataOut[3427]),
.io_parallelOut_3428(dataOut[3428]),
.io_parallelOut_3429(dataOut[3429]),
.io_parallelOut_3430(dataOut[3430]),
.io_parallelOut_3431(dataOut[3431]),
.io_parallelOut_3432(dataOut[3432]),
.io_parallelOut_3433(dataOut[3433]),
.io_parallelOut_3434(dataOut[3434]),
.io_parallelOut_3435(dataOut[3435]),
.io_parallelOut_3436(dataOut[3436]),
.io_parallelOut_3437(dataOut[3437]),
.io_parallelOut_3438(dataOut[3438]),
.io_parallelOut_3439(dataOut[3439]),
.io_parallelOut_3440(dataOut[3440]),
.io_parallelOut_3441(dataOut[3441]),
.io_parallelOut_3442(dataOut[3442]),
.io_parallelOut_3443(dataOut[3443]),
.io_parallelOut_3444(dataOut[3444]),
.io_parallelOut_3445(dataOut[3445]),
.io_parallelOut_3446(dataOut[3446]),
.io_parallelOut_3447(dataOut[3447]),
.io_parallelOut_3448(dataOut[3448]),
.io_parallelOut_3449(dataOut[3449]),
.io_parallelOut_3450(dataOut[3450]),
.io_parallelOut_3451(dataOut[3451]),
.io_parallelOut_3452(dataOut[3452]),
.io_parallelOut_3453(dataOut[3453]),
.io_parallelOut_3454(dataOut[3454]),
.io_parallelOut_3455(dataOut[3455]),
.io_parallelOut_3456(dataOut[3456]),
.io_parallelOut_3457(dataOut[3457]),
.io_parallelOut_3458(dataOut[3458]),
.io_parallelOut_3459(dataOut[3459]),
.io_parallelOut_3460(dataOut[3460]),
.io_parallelOut_3461(dataOut[3461]),
.io_parallelOut_3462(dataOut[3462]),
.io_parallelOut_3463(dataOut[3463]),
.io_parallelOut_3464(dataOut[3464]),
.io_parallelOut_3465(dataOut[3465]),
.io_parallelOut_3466(dataOut[3466]),
.io_parallelOut_3467(dataOut[3467]),
.io_parallelOut_3468(dataOut[3468]),
.io_parallelOut_3469(dataOut[3469]),
.io_parallelOut_3470(dataOut[3470]),
.io_parallelOut_3471(dataOut[3471]),
.io_parallelOut_3472(dataOut[3472]),
.io_parallelOut_3473(dataOut[3473]),
.io_parallelOut_3474(dataOut[3474]),
.io_parallelOut_3475(dataOut[3475]),
.io_parallelOut_3476(dataOut[3476]),
.io_parallelOut_3477(dataOut[3477]),
.io_parallelOut_3478(dataOut[3478]),
.io_parallelOut_3479(dataOut[3479]),
.io_parallelOut_3480(dataOut[3480]),
.io_parallelOut_3481(dataOut[3481]),
.io_parallelOut_3482(dataOut[3482]),
.io_parallelOut_3483(dataOut[3483]),
.io_parallelOut_3484(dataOut[3484]),
.io_parallelOut_3485(dataOut[3485]),
.io_parallelOut_3486(dataOut[3486]),
.io_parallelOut_3487(dataOut[3487]),
.io_parallelOut_3488(dataOut[3488]),
.io_parallelOut_3489(dataOut[3489]),
.io_parallelOut_3490(dataOut[3490]),
.io_parallelOut_3491(dataOut[3491]),
.io_parallelOut_3492(dataOut[3492]),
.io_parallelOut_3493(dataOut[3493]),
.io_parallelOut_3494(dataOut[3494]),
.io_parallelOut_3495(dataOut[3495]),
.io_parallelOut_3496(dataOut[3496]),
.io_parallelOut_3497(dataOut[3497]),
.io_parallelOut_3498(dataOut[3498]),
.io_parallelOut_3499(dataOut[3499]),
.io_parallelOut_3500(dataOut[3500]),
.io_parallelOut_3501(dataOut[3501]),
.io_parallelOut_3502(dataOut[3502]),
.io_parallelOut_3503(dataOut[3503]),
.io_parallelOut_3504(dataOut[3504]),
.io_parallelOut_3505(dataOut[3505]),
.io_parallelOut_3506(dataOut[3506]),
.io_parallelOut_3507(dataOut[3507]),
.io_parallelOut_3508(dataOut[3508]),
.io_parallelOut_3509(dataOut[3509]),
.io_parallelOut_3510(dataOut[3510]),
.io_parallelOut_3511(dataOut[3511]),
.io_parallelOut_3512(dataOut[3512]),
.io_parallelOut_3513(dataOut[3513]),
.io_parallelOut_3514(dataOut[3514]),
.io_parallelOut_3515(dataOut[3515]),
.io_parallelOut_3516(dataOut[3516]),
.io_parallelOut_3517(dataOut[3517]),
.io_parallelOut_3518(dataOut[3518]),
.io_parallelOut_3519(dataOut[3519]),
.io_parallelOut_3520(dataOut[3520]),
.io_parallelOut_3521(dataOut[3521]),
.io_parallelOut_3522(dataOut[3522]),
.io_parallelOut_3523(dataOut[3523]),
.io_parallelOut_3524(dataOut[3524]),
.io_parallelOut_3525(dataOut[3525]),
.io_parallelOut_3526(dataOut[3526]),
.io_parallelOut_3527(dataOut[3527]),
.io_parallelOut_3528(dataOut[3528]),
.io_parallelOut_3529(dataOut[3529]),
.io_parallelOut_3530(dataOut[3530]),
.io_parallelOut_3531(dataOut[3531]),
.io_parallelOut_3532(dataOut[3532]),
.io_parallelOut_3533(dataOut[3533]),
.io_parallelOut_3534(dataOut[3534]),
.io_parallelOut_3535(dataOut[3535]),
.io_parallelOut_3536(dataOut[3536]),
.io_parallelOut_3537(dataOut[3537]),
.io_parallelOut_3538(dataOut[3538]),
.io_parallelOut_3539(dataOut[3539]),
.io_parallelOut_3540(dataOut[3540]),
.io_parallelOut_3541(dataOut[3541]),
.io_parallelOut_3542(dataOut[3542]),
.io_parallelOut_3543(dataOut[3543]),
.io_parallelOut_3544(dataOut[3544]),
.io_parallelOut_3545(dataOut[3545]),
.io_parallelOut_3546(dataOut[3546]),
.io_parallelOut_3547(dataOut[3547]),
.io_parallelOut_3548(dataOut[3548]),
.io_parallelOut_3549(dataOut[3549]),
.io_parallelOut_3550(dataOut[3550]),
.io_parallelOut_3551(dataOut[3551]),
.io_parallelOut_3552(dataOut[3552]),
.io_parallelOut_3553(dataOut[3553]),
.io_parallelOut_3554(dataOut[3554]),
.io_parallelOut_3555(dataOut[3555]),
.io_parallelOut_3556(dataOut[3556]),
.io_parallelOut_3557(dataOut[3557]),
.io_parallelOut_3558(dataOut[3558]),
.io_parallelOut_3559(dataOut[3559]),
.io_parallelOut_3560(dataOut[3560]),
.io_parallelOut_3561(dataOut[3561]),
.io_parallelOut_3562(dataOut[3562]),
.io_parallelOut_3563(dataOut[3563]),
.io_parallelOut_3564(dataOut[3564]),
.io_parallelOut_3565(dataOut[3565]),
.io_parallelOut_3566(dataOut[3566]),
.io_parallelOut_3567(dataOut[3567]),
.io_parallelOut_3568(dataOut[3568]),
.io_parallelOut_3569(dataOut[3569]),
.io_parallelOut_3570(dataOut[3570]),
.io_parallelOut_3571(dataOut[3571]),
.io_parallelOut_3572(dataOut[3572]),
.io_parallelOut_3573(dataOut[3573]),
.io_parallelOut_3574(dataOut[3574]),
.io_parallelOut_3575(dataOut[3575]),
.io_parallelOut_3576(dataOut[3576]),
.io_parallelOut_3577(dataOut[3577]),
.io_parallelOut_3578(dataOut[3578]),
.io_parallelOut_3579(dataOut[3579]),
.io_parallelOut_3580(dataOut[3580]),
.io_parallelOut_3581(dataOut[3581]),
.io_parallelOut_3582(dataOut[3582]),
.io_parallelOut_3583(dataOut[3583]),
.io_parallelOut_3584(dataOut[3584]),
.io_parallelOut_3585(dataOut[3585]),
.io_parallelOut_3586(dataOut[3586]),
.io_parallelOut_3587(dataOut[3587]),
.io_parallelOut_3588(dataOut[3588]),
.io_parallelOut_3589(dataOut[3589]),
.io_parallelOut_3590(dataOut[3590]),
.io_parallelOut_3591(dataOut[3591]),
.io_parallelOut_3592(dataOut[3592]),
.io_parallelOut_3593(dataOut[3593]),
.io_parallelOut_3594(dataOut[3594]),
.io_parallelOut_3595(dataOut[3595]),
.io_parallelOut_3596(dataOut[3596]),
.io_parallelOut_3597(dataOut[3597]),
.io_parallelOut_3598(dataOut[3598]),
.io_parallelOut_3599(dataOut[3599]),
.io_parallelOut_3600(dataOut[3600]),
.io_parallelOut_3601(dataOut[3601]),
.io_parallelOut_3602(dataOut[3602]),
.io_parallelOut_3603(dataOut[3603]),
.io_parallelOut_3604(dataOut[3604]),
.io_parallelOut_3605(dataOut[3605]),
.io_parallelOut_3606(dataOut[3606]),
.io_parallelOut_3607(dataOut[3607]),
.io_parallelOut_3608(dataOut[3608]),
.io_parallelOut_3609(dataOut[3609]),
.io_parallelOut_3610(dataOut[3610]),
.io_parallelOut_3611(dataOut[3611]),
.io_parallelOut_3612(dataOut[3612]),
.io_parallelOut_3613(dataOut[3613]),
.io_parallelOut_3614(dataOut[3614]),
.io_parallelOut_3615(dataOut[3615]),
.io_parallelOut_3616(dataOut[3616]),
.io_parallelOut_3617(dataOut[3617]),
.io_parallelOut_3618(dataOut[3618]),
.io_parallelOut_3619(dataOut[3619]),
.io_parallelOut_3620(dataOut[3620]),
.io_parallelOut_3621(dataOut[3621]),
.io_parallelOut_3622(dataOut[3622]),
.io_parallelOut_3623(dataOut[3623]),
.io_parallelOut_3624(dataOut[3624]),
.io_parallelOut_3625(dataOut[3625]),
.io_parallelOut_3626(dataOut[3626]),
.io_parallelOut_3627(dataOut[3627]),
.io_parallelOut_3628(dataOut[3628]),
.io_parallelOut_3629(dataOut[3629]),
.io_parallelOut_3630(dataOut[3630]),
.io_parallelOut_3631(dataOut[3631]),
.io_parallelOut_3632(dataOut[3632]),
.io_parallelOut_3633(dataOut[3633]),
.io_parallelOut_3634(dataOut[3634]),
.io_parallelOut_3635(dataOut[3635]),
.io_parallelOut_3636(dataOut[3636]),
.io_parallelOut_3637(dataOut[3637]),
.io_parallelOut_3638(dataOut[3638]),
.io_parallelOut_3639(dataOut[3639]),
.io_parallelOut_3640(dataOut[3640]),
.io_parallelOut_3641(dataOut[3641]),
.io_parallelOut_3642(dataOut[3642]),
.io_parallelOut_3643(dataOut[3643]),
.io_parallelOut_3644(dataOut[3644]),
.io_parallelOut_3645(dataOut[3645]),
.io_parallelOut_3646(dataOut[3646]),
.io_parallelOut_3647(dataOut[3647]),
.io_parallelOut_3648(dataOut[3648]),
.io_parallelOut_3649(dataOut[3649]),
.io_parallelOut_3650(dataOut[3650]),
.io_parallelOut_3651(dataOut[3651]),
.io_parallelOut_3652(dataOut[3652]),
.io_parallelOut_3653(dataOut[3653]),
.io_parallelOut_3654(dataOut[3654]),
.io_parallelOut_3655(dataOut[3655]),
.io_parallelOut_3656(dataOut[3656]),
.io_parallelOut_3657(dataOut[3657]),
.io_parallelOut_3658(dataOut[3658]),
.io_parallelOut_3659(dataOut[3659]),
.io_parallelOut_3660(dataOut[3660]),
.io_parallelOut_3661(dataOut[3661]),
.io_parallelOut_3662(dataOut[3662]),
.io_parallelOut_3663(dataOut[3663]),
.io_parallelOut_3664(dataOut[3664]),
.io_parallelOut_3665(dataOut[3665]),
.io_parallelOut_3666(dataOut[3666]),
.io_parallelOut_3667(dataOut[3667]),
.io_parallelOut_3668(dataOut[3668]),
.io_parallelOut_3669(dataOut[3669]),
.io_parallelOut_3670(dataOut[3670]),
.io_parallelOut_3671(dataOut[3671]),
.io_parallelOut_3672(dataOut[3672]),
.io_parallelOut_3673(dataOut[3673]),
.io_parallelOut_3674(dataOut[3674]),
.io_parallelOut_3675(dataOut[3675]),
.io_parallelOut_3676(dataOut[3676]),
.io_parallelOut_3677(dataOut[3677]),
.io_parallelOut_3678(dataOut[3678]),
.io_parallelOut_3679(dataOut[3679]),
.io_parallelOut_3680(dataOut[3680]),
.io_parallelOut_3681(dataOut[3681]),
.io_parallelOut_3682(dataOut[3682]),
.io_parallelOut_3683(dataOut[3683]),
.io_parallelOut_3684(dataOut[3684]),
.io_parallelOut_3685(dataOut[3685]),
.io_parallelOut_3686(dataOut[3686]),
.io_parallelOut_3687(dataOut[3687]),
.io_parallelOut_3688(dataOut[3688]),
.io_parallelOut_3689(dataOut[3689]),
.io_parallelOut_3690(dataOut[3690]),
.io_parallelOut_3691(dataOut[3691]),
.io_parallelOut_3692(dataOut[3692]),
.io_parallelOut_3693(dataOut[3693]),
.io_parallelOut_3694(dataOut[3694]),
.io_parallelOut_3695(dataOut[3695]),
.io_parallelOut_3696(dataOut[3696]),
.io_parallelOut_3697(dataOut[3697]),
.io_parallelOut_3698(dataOut[3698]),
.io_parallelOut_3699(dataOut[3699]),
.io_parallelOut_3700(dataOut[3700]),
.io_parallelOut_3701(dataOut[3701]),
.io_parallelOut_3702(dataOut[3702]),
.io_parallelOut_3703(dataOut[3703]),
.io_parallelOut_3704(dataOut[3704]),
.io_parallelOut_3705(dataOut[3705]),
.io_parallelOut_3706(dataOut[3706]),
.io_parallelOut_3707(dataOut[3707]),
.io_parallelOut_3708(dataOut[3708]),
.io_parallelOut_3709(dataOut[3709]),
.io_parallelOut_3710(dataOut[3710]),
.io_parallelOut_3711(dataOut[3711]),
.io_parallelOut_3712(dataOut[3712]),
.io_parallelOut_3713(dataOut[3713]),
.io_parallelOut_3714(dataOut[3714]),
.io_parallelOut_3715(dataOut[3715]),
.io_parallelOut_3716(dataOut[3716]),
.io_parallelOut_3717(dataOut[3717]),
.io_parallelOut_3718(dataOut[3718]),
.io_parallelOut_3719(dataOut[3719]),
.io_parallelOut_3720(dataOut[3720]),
.io_parallelOut_3721(dataOut[3721]),
.io_parallelOut_3722(dataOut[3722]),
.io_parallelOut_3723(dataOut[3723]),
.io_parallelOut_3724(dataOut[3724]),
.io_parallelOut_3725(dataOut[3725]),
.io_parallelOut_3726(dataOut[3726]),
.io_parallelOut_3727(dataOut[3727]),
.io_parallelOut_3728(dataOut[3728]),
.io_parallelOut_3729(dataOut[3729]),
.io_parallelOut_3730(dataOut[3730]),
.io_parallelOut_3731(dataOut[3731]),
.io_parallelOut_3732(dataOut[3732]),
.io_parallelOut_3733(dataOut[3733]),
.io_parallelOut_3734(dataOut[3734]),
.io_parallelOut_3735(dataOut[3735]),
.io_parallelOut_3736(dataOut[3736]),
.io_parallelOut_3737(dataOut[3737]),
.io_parallelOut_3738(dataOut[3738]),
.io_parallelOut_3739(dataOut[3739]),
.io_parallelOut_3740(dataOut[3740]),
.io_parallelOut_3741(dataOut[3741]),
.io_parallelOut_3742(dataOut[3742]),
.io_parallelOut_3743(dataOut[3743]),
.io_parallelOut_3744(dataOut[3744]),
.io_parallelOut_3745(dataOut[3745]),
.io_parallelOut_3746(dataOut[3746]),
.io_parallelOut_3747(dataOut[3747]),
.io_parallelOut_3748(dataOut[3748]),
.io_parallelOut_3749(dataOut[3749]),
.io_parallelOut_3750(dataOut[3750]),
.io_parallelOut_3751(dataOut[3751]),
.io_parallelOut_3752(dataOut[3752]),
.io_parallelOut_3753(dataOut[3753]),
.io_parallelOut_3754(dataOut[3754]),
.io_parallelOut_3755(dataOut[3755]),
.io_parallelOut_3756(dataOut[3756]),
.io_parallelOut_3757(dataOut[3757]),
.io_parallelOut_3758(dataOut[3758]),
.io_parallelOut_3759(dataOut[3759]),
.io_parallelOut_3760(dataOut[3760]),
.io_parallelOut_3761(dataOut[3761]),
.io_parallelOut_3762(dataOut[3762]),
.io_parallelOut_3763(dataOut[3763]),
.io_parallelOut_3764(dataOut[3764]),
.io_parallelOut_3765(dataOut[3765]),
.io_parallelOut_3766(dataOut[3766]),
.io_parallelOut_3767(dataOut[3767]),
.io_parallelOut_3768(dataOut[3768]),
.io_parallelOut_3769(dataOut[3769]),
.io_parallelOut_3770(dataOut[3770]),
.io_parallelOut_3771(dataOut[3771]),
.io_parallelOut_3772(dataOut[3772]),
.io_parallelOut_3773(dataOut[3773]),
.io_parallelOut_3774(dataOut[3774]),
.io_parallelOut_3775(dataOut[3775]),
.io_parallelOut_3776(dataOut[3776]),
.io_parallelOut_3777(dataOut[3777]),
.io_parallelOut_3778(dataOut[3778]),
.io_parallelOut_3779(dataOut[3779]),
.io_parallelOut_3780(dataOut[3780]),
.io_parallelOut_3781(dataOut[3781]),
.io_parallelOut_3782(dataOut[3782]),
.io_parallelOut_3783(dataOut[3783]),
.io_parallelOut_3784(dataOut[3784]),
.io_parallelOut_3785(dataOut[3785]),
.io_parallelOut_3786(dataOut[3786]),
.io_parallelOut_3787(dataOut[3787]),
.io_parallelOut_3788(dataOut[3788]),
.io_parallelOut_3789(dataOut[3789]),
.io_parallelOut_3790(dataOut[3790]),
.io_parallelOut_3791(dataOut[3791]),
.io_parallelOut_3792(dataOut[3792]),
.io_parallelOut_3793(dataOut[3793]),
.io_parallelOut_3794(dataOut[3794]),
.io_parallelOut_3795(dataOut[3795]),
.io_parallelOut_3796(dataOut[3796]),
.io_parallelOut_3797(dataOut[3797]),
.io_parallelOut_3798(dataOut[3798]),
.io_parallelOut_3799(dataOut[3799]),
.io_parallelOut_3800(dataOut[3800]),
.io_parallelOut_3801(dataOut[3801]),
.io_parallelOut_3802(dataOut[3802]),
.io_parallelOut_3803(dataOut[3803]),
.io_parallelOut_3804(dataOut[3804]),
.io_parallelOut_3805(dataOut[3805]),
.io_parallelOut_3806(dataOut[3806]),
.io_parallelOut_3807(dataOut[3807]),
.io_parallelOut_3808(dataOut[3808]),
.io_parallelOut_3809(dataOut[3809]),
.io_parallelOut_3810(dataOut[3810]),
.io_parallelOut_3811(dataOut[3811]),
.io_parallelOut_3812(dataOut[3812]),
.io_parallelOut_3813(dataOut[3813]),
.io_parallelOut_3814(dataOut[3814]),
.io_parallelOut_3815(dataOut[3815]),
.io_parallelOut_3816(dataOut[3816]),
.io_parallelOut_3817(dataOut[3817]),
.io_parallelOut_3818(dataOut[3818]),
.io_parallelOut_3819(dataOut[3819]),
.io_parallelOut_3820(dataOut[3820]),
.io_parallelOut_3821(dataOut[3821]),
.io_parallelOut_3822(dataOut[3822]),
.io_parallelOut_3823(dataOut[3823]),
.io_parallelOut_3824(dataOut[3824]),
.io_parallelOut_3825(dataOut[3825]),
.io_parallelOut_3826(dataOut[3826]),
.io_parallelOut_3827(dataOut[3827]),
.io_parallelOut_3828(dataOut[3828]),
.io_parallelOut_3829(dataOut[3829]),
.io_parallelOut_3830(dataOut[3830]),
.io_parallelOut_3831(dataOut[3831]),
.io_parallelOut_3832(dataOut[3832]),
.io_parallelOut_3833(dataOut[3833]),
.io_parallelOut_3834(dataOut[3834]),
.io_parallelOut_3835(dataOut[3835]),
.io_parallelOut_3836(dataOut[3836]),
.io_parallelOut_3837(dataOut[3837]),
.io_parallelOut_3838(dataOut[3838]),
.io_parallelOut_3839(dataOut[3839]),
.io_parallelOut_3840(dataOut[3840]),
.io_parallelOut_3841(dataOut[3841]),
.io_parallelOut_3842(dataOut[3842]),
.io_parallelOut_3843(dataOut[3843]),
.io_parallelOut_3844(dataOut[3844]),
.io_parallelOut_3845(dataOut[3845]),
.io_parallelOut_3846(dataOut[3846]),
.io_parallelOut_3847(dataOut[3847]),
.io_parallelOut_3848(dataOut[3848]),
.io_parallelOut_3849(dataOut[3849]),
.io_parallelOut_3850(dataOut[3850]),
.io_parallelOut_3851(dataOut[3851]),
.io_parallelOut_3852(dataOut[3852]),
.io_parallelOut_3853(dataOut[3853]),
.io_parallelOut_3854(dataOut[3854]),
.io_parallelOut_3855(dataOut[3855]),
.io_parallelOut_3856(dataOut[3856]),
.io_parallelOut_3857(dataOut[3857]),
.io_parallelOut_3858(dataOut[3858]),
.io_parallelOut_3859(dataOut[3859]),
.io_parallelOut_3860(dataOut[3860]),
.io_parallelOut_3861(dataOut[3861]),
.io_parallelOut_3862(dataOut[3862]),
.io_parallelOut_3863(dataOut[3863]),
.io_parallelOut_3864(dataOut[3864]),
.io_parallelOut_3865(dataOut[3865]),
.io_parallelOut_3866(dataOut[3866]),
.io_parallelOut_3867(dataOut[3867]),
.io_parallelOut_3868(dataOut[3868]),
.io_parallelOut_3869(dataOut[3869]),
.io_parallelOut_3870(dataOut[3870]),
.io_parallelOut_3871(dataOut[3871]),
.io_parallelOut_3872(dataOut[3872]),
.io_parallelOut_3873(dataOut[3873]),
.io_parallelOut_3874(dataOut[3874]),
.io_parallelOut_3875(dataOut[3875]),
.io_parallelOut_3876(dataOut[3876]),
.io_parallelOut_3877(dataOut[3877]),
.io_parallelOut_3878(dataOut[3878]),
.io_parallelOut_3879(dataOut[3879]),
.io_parallelOut_3880(dataOut[3880]),
.io_parallelOut_3881(dataOut[3881]),
.io_parallelOut_3882(dataOut[3882]),
.io_parallelOut_3883(dataOut[3883]),
.io_parallelOut_3884(dataOut[3884]),
.io_parallelOut_3885(dataOut[3885]),
.io_parallelOut_3886(dataOut[3886]),
.io_parallelOut_3887(dataOut[3887]),
.io_parallelOut_3888(dataOut[3888]),
.io_parallelOut_3889(dataOut[3889]),
.io_parallelOut_3890(dataOut[3890]),
.io_parallelOut_3891(dataOut[3891]),
.io_parallelOut_3892(dataOut[3892]),
.io_parallelOut_3893(dataOut[3893]),
.io_parallelOut_3894(dataOut[3894]),
.io_parallelOut_3895(dataOut[3895]),
.io_parallelOut_3896(dataOut[3896]),
.io_parallelOut_3897(dataOut[3897]),
.io_parallelOut_3898(dataOut[3898]),
.io_parallelOut_3899(dataOut[3899]),
.io_parallelOut_3900(dataOut[3900]),
.io_parallelOut_3901(dataOut[3901]),
.io_parallelOut_3902(dataOut[3902]),
.io_parallelOut_3903(dataOut[3903]),
.io_parallelOut_3904(dataOut[3904]),
.io_parallelOut_3905(dataOut[3905]),
.io_parallelOut_3906(dataOut[3906]),
.io_parallelOut_3907(dataOut[3907]),
.io_parallelOut_3908(dataOut[3908]),
.io_parallelOut_3909(dataOut[3909]),
.io_parallelOut_3910(dataOut[3910]),
.io_parallelOut_3911(dataOut[3911]),
.io_parallelOut_3912(dataOut[3912]),
.io_parallelOut_3913(dataOut[3913]),
.io_parallelOut_3914(dataOut[3914]),
.io_parallelOut_3915(dataOut[3915]),
.io_parallelOut_3916(dataOut[3916]),
.io_parallelOut_3917(dataOut[3917]),
.io_parallelOut_3918(dataOut[3918]),
.io_parallelOut_3919(dataOut[3919]),
.io_parallelOut_3920(dataOut[3920]),
.io_parallelOut_3921(dataOut[3921]),
.io_parallelOut_3922(dataOut[3922]),
.io_parallelOut_3923(dataOut[3923]),
.io_parallelOut_3924(dataOut[3924]),
.io_parallelOut_3925(dataOut[3925]),
.io_parallelOut_3926(dataOut[3926]),
.io_parallelOut_3927(dataOut[3927]),
.io_parallelOut_3928(dataOut[3928]),
.io_parallelOut_3929(dataOut[3929]),
.io_parallelOut_3930(dataOut[3930]),
.io_parallelOut_3931(dataOut[3931]),
.io_parallelOut_3932(dataOut[3932]),
.io_parallelOut_3933(dataOut[3933]),
.io_parallelOut_3934(dataOut[3934]),
.io_parallelOut_3935(dataOut[3935]),
.io_parallelOut_3936(dataOut[3936]),
.io_parallelOut_3937(dataOut[3937]),
.io_parallelOut_3938(dataOut[3938]),
.io_parallelOut_3939(dataOut[3939]),
.io_parallelOut_3940(dataOut[3940]),
.io_parallelOut_3941(dataOut[3941]),
.io_parallelOut_3942(dataOut[3942]),
.io_parallelOut_3943(dataOut[3943]),
.io_parallelOut_3944(dataOut[3944]),
.io_parallelOut_3945(dataOut[3945]),
.io_parallelOut_3946(dataOut[3946]),
.io_parallelOut_3947(dataOut[3947]),
.io_parallelOut_3948(dataOut[3948]),
.io_parallelOut_3949(dataOut[3949]),
.io_parallelOut_3950(dataOut[3950]),
.io_parallelOut_3951(dataOut[3951]),
.io_parallelOut_3952(dataOut[3952]),
.io_parallelOut_3953(dataOut[3953]),
.io_parallelOut_3954(dataOut[3954]),
.io_parallelOut_3955(dataOut[3955]),
.io_parallelOut_3956(dataOut[3956]),
.io_parallelOut_3957(dataOut[3957]),
.io_parallelOut_3958(dataOut[3958]),
.io_parallelOut_3959(dataOut[3959]),
.io_parallelOut_3960(dataOut[3960]),
.io_parallelOut_3961(dataOut[3961]),
.io_parallelOut_3962(dataOut[3962]),
.io_parallelOut_3963(dataOut[3963]),
.io_parallelOut_3964(dataOut[3964]),
.io_parallelOut_3965(dataOut[3965]),
.io_parallelOut_3966(dataOut[3966]),
.io_parallelOut_3967(dataOut[3967]),
.io_parallelOut_3968(dataOut[3968]),
.io_parallelOut_3969(dataOut[3969]),
.io_parallelOut_3970(dataOut[3970]),
.io_parallelOut_3971(dataOut[3971]),
.io_parallelOut_3972(dataOut[3972]),
.io_parallelOut_3973(dataOut[3973]),
.io_parallelOut_3974(dataOut[3974]),
.io_parallelOut_3975(dataOut[3975]),
.io_parallelOut_3976(dataOut[3976]),
.io_parallelOut_3977(dataOut[3977]),
.io_parallelOut_3978(dataOut[3978]),
.io_parallelOut_3979(dataOut[3979]),
.io_parallelOut_3980(dataOut[3980]),
.io_parallelOut_3981(dataOut[3981]),
.io_parallelOut_3982(dataOut[3982]),
.io_parallelOut_3983(dataOut[3983]),
.io_parallelOut_3984(dataOut[3984]),
.io_parallelOut_3985(dataOut[3985]),
.io_parallelOut_3986(dataOut[3986]),
.io_parallelOut_3987(dataOut[3987]),
.io_parallelOut_3988(dataOut[3988]),
.io_parallelOut_3989(dataOut[3989]),
.io_parallelOut_3990(dataOut[3990]),
.io_parallelOut_3991(dataOut[3991]),
.io_parallelOut_3992(dataOut[3992]),
.io_parallelOut_3993(dataOut[3993]),
.io_parallelOut_3994(dataOut[3994]),
.io_parallelOut_3995(dataOut[3995]),
.io_parallelOut_3996(dataOut[3996]),
.io_parallelOut_3997(dataOut[3997]),
.io_parallelOut_3998(dataOut[3998]),
.io_parallelOut_3999(dataOut[3999]),
.io_parallelOut_4000(dataOut[4000]),
.io_parallelOut_4001(dataOut[4001]),
.io_parallelOut_4002(dataOut[4002]),
.io_parallelOut_4003(dataOut[4003]),
.io_parallelOut_4004(dataOut[4004]),
.io_parallelOut_4005(dataOut[4005]),
.io_parallelOut_4006(dataOut[4006]),
.io_parallelOut_4007(dataOut[4007]),
.io_parallelOut_4008(dataOut[4008]),
.io_parallelOut_4009(dataOut[4009]),
.io_parallelOut_4010(dataOut[4010]),
.io_parallelOut_4011(dataOut[4011]),
.io_parallelOut_4012(dataOut[4012]),
.io_parallelOut_4013(dataOut[4013]),
.io_parallelOut_4014(dataOut[4014]),
.io_parallelOut_4015(dataOut[4015]),
.io_parallelOut_4016(dataOut[4016]),
.io_parallelOut_4017(dataOut[4017]),
.io_parallelOut_4018(dataOut[4018]),
.io_parallelOut_4019(dataOut[4019]),
.io_parallelOut_4020(dataOut[4020]),
.io_parallelOut_4021(dataOut[4021]),
.io_parallelOut_4022(dataOut[4022]),
.io_parallelOut_4023(dataOut[4023]),
.io_parallelOut_4024(dataOut[4024]),
.io_parallelOut_4025(dataOut[4025]),
.io_parallelOut_4026(dataOut[4026]),
.io_parallelOut_4027(dataOut[4027]),
.io_parallelOut_4028(dataOut[4028]),
.io_parallelOut_4029(dataOut[4029]),
.io_parallelOut_4030(dataOut[4030]),
.io_parallelOut_4031(dataOut[4031]),
.io_parallelOut_4032(dataOut[4032]),
.io_parallelOut_4033(dataOut[4033]),
.io_parallelOut_4034(dataOut[4034]),
.io_parallelOut_4035(dataOut[4035]),
.io_parallelOut_4036(dataOut[4036]),
.io_parallelOut_4037(dataOut[4037]),
.io_parallelOut_4038(dataOut[4038]),
.io_parallelOut_4039(dataOut[4039]),
.io_parallelOut_4040(dataOut[4040]),
.io_parallelOut_4041(dataOut[4041]),
.io_parallelOut_4042(dataOut[4042]),
.io_parallelOut_4043(dataOut[4043]),
.io_parallelOut_4044(dataOut[4044]),
.io_parallelOut_4045(dataOut[4045]),
.io_parallelOut_4046(dataOut[4046]),
.io_parallelOut_4047(dataOut[4047]),
.io_parallelOut_4048(dataOut[4048]),
.io_parallelOut_4049(dataOut[4049]),
.io_parallelOut_4050(dataOut[4050]),
.io_parallelOut_4051(dataOut[4051]),
.io_parallelOut_4052(dataOut[4052]),
.io_parallelOut_4053(dataOut[4053]),
.io_parallelOut_4054(dataOut[4054]),
.io_parallelOut_4055(dataOut[4055]),
.io_parallelOut_4056(dataOut[4056]),
.io_parallelOut_4057(dataOut[4057]),
.io_parallelOut_4058(dataOut[4058]),
.io_parallelOut_4059(dataOut[4059]),
.io_parallelOut_4060(dataOut[4060]),
.io_parallelOut_4061(dataOut[4061]),
.io_parallelOut_4062(dataOut[4062]),
.io_parallelOut_4063(dataOut[4063]),
.io_parallelOut_4064(dataOut[4064]),
.io_parallelOut_4065(dataOut[4065]),
.io_parallelOut_4066(dataOut[4066]),
.io_parallelOut_4067(dataOut[4067]),
.io_parallelOut_4068(dataOut[4068]),
.io_parallelOut_4069(dataOut[4069]),
.io_parallelOut_4070(dataOut[4070]),
.io_parallelOut_4071(dataOut[4071]),
.io_parallelOut_4072(dataOut[4072]),
.io_parallelOut_4073(dataOut[4073]),
.io_parallelOut_4074(dataOut[4074]),
.io_parallelOut_4075(dataOut[4075]),
.io_parallelOut_4076(dataOut[4076]),
.io_parallelOut_4077(dataOut[4077]),
.io_parallelOut_4078(dataOut[4078]),
.io_parallelOut_4079(dataOut[4079]),
.io_parallelOut_4080(dataOut[4080]),
.io_parallelOut_4081(dataOut[4081]),
.io_parallelOut_4082(dataOut[4082]),
.io_parallelOut_4083(dataOut[4083]),
.io_parallelOut_4084(dataOut[4084]),
.io_parallelOut_4085(dataOut[4085]),
.io_parallelOut_4086(dataOut[4086]),
.io_parallelOut_4087(dataOut[4087]),
.io_parallelOut_4088(dataOut[4088]),
.io_parallelOut_4089(dataOut[4089]),
.io_parallelOut_4090(dataOut[4090]),
.io_parallelOut_4091(dataOut[4091]),
.io_parallelOut_4092(dataOut[4092]),
.io_parallelOut_4093(dataOut[4093]),
.io_parallelOut_4094(dataOut[4094]),
.io_parallelOut_4095(dataOut[4095]),
.io_matchBytes_0(matchBytes[0]),
.io_matchBytes_1(matchBytes[1]),
.io_matchBytes_2(matchBytes[2]),
.io_matchBytes_3(matchBytes[3]),
.io_matchBytes_4(matchBytes[4]),
.io_matchBytes_5(matchBytes[5]),
.io_matchBytes_6(matchBytes[6]),
.io_matchBytes_7(matchBytes[7]),
.io_matchBytes_8(matchBytes[8]),
.io_matchBytes_9(matchBytes[9]),
.io_matchBytes_10(matchBytes[10]),
.io_matchBytes_11(matchBytes[11]),
.io_matchBytes_12(matchBytes[12]),
.io_matchBytes_13(matchBytes[13]),
.io_matchBytes_14(matchBytes[14]),
.io_matchBytes_15(matchBytes[15]),
.io_matchBytes_16(matchBytes[16]),
.io_matchBytes_17(matchBytes[17]),
.io_matchBytes_18(matchBytes[18]),
.io_matchBytes_19(matchBytes[19]),
.io_matchBytes_20(matchBytes[20]),
.io_matchBytes_21(matchBytes[21]),
.io_matchBytes_22(matchBytes[22]),
.io_matchBytes_23(matchBytes[23]),
.io_matchBytes_24(matchBytes[24]),
.io_matchBytes_25(matchBytes[25]),
.io_matchBytes_26(matchBytes[26]),
.io_matchBytes_27(matchBytes[27]),
.io_matchBytes_28(matchBytes[28]),
.io_matchBytes_29(matchBytes[29]),
.io_matchBytes_30(matchBytes[30]),
.io_matchBytes_31(matchBytes[31]),
.io_matchBytes_32(matchBytes[32]),
.io_matchBytes_33(matchBytes[33]),
.io_matchBytes_34(matchBytes[34]),
.io_matchBytes_35(matchBytes[35]),
.io_matchBytes_36(matchBytes[36]),
.io_matchBytes_37(matchBytes[37]),
.io_matchBytes_38(matchBytes[38]),
.io_matchBytes_39(matchBytes[39]),
.io_matchBytes_40(matchBytes[40]),
.io_matchBytes_41(matchBytes[41]),
.io_matchBytes_42(matchBytes[42]),
.io_matchBytes_43(matchBytes[43]),
.io_matchBytes_44(matchBytes[44]),
.io_matchBytes_45(matchBytes[45]),
.io_matchBytes_46(matchBytes[46]),
.io_matchBytes_47(matchBytes[47]),
.io_matchBytes_48(matchBytes[48]),
.io_matchBytes_49(matchBytes[49]),
.io_matchBytes_50(matchBytes[50]),
.io_matchBytes_51(matchBytes[51]),
.io_matchBytes_52(matchBytes[52]),
.io_matchBytes_53(matchBytes[53]),
.io_matchBytes_54(matchBytes[54]),
.io_matchBytes_55(matchBytes[55]),
.io_matchBytes_56(matchBytes[56]),
.io_matchBytes_57(matchBytes[57]),
.io_matchBytes_58(matchBytes[58]),
.io_matchBytes_59(matchBytes[59]),
.io_matchBytes_60(matchBytes[60]),
.io_matchBytes_61(matchBytes[61]),
.io_matchBytes_62(matchBytes[62]),
.io_matchBytes_63(matchBytes[63]),
.io_matchBytes_64(matchBytes[64]),
.io_matchBytes_65(matchBytes[65]),
.io_matchBytes_66(matchBytes[66]),
.io_matchBytes_67(matchBytes[67]),
.io_matchBytes_68(matchBytes[68]),
.io_matchBytes_69(matchBytes[69]),
.io_matchBytes_70(matchBytes[70]),
.io_matchBytes_71(matchBytes[71]),
.io_matchBytes_72(matchBytes[72]),
.io_matchBytes_73(matchBytes[73]),
.io_matchBytes_74(matchBytes[74]),
.io_matchBytes_75(matchBytes[75]),
.io_matchBytes_76(matchBytes[76]),
.io_matchBytes_77(matchBytes[77]),
.io_matchBytes_78(matchBytes[78]),
.io_matchBytes_79(matchBytes[79]),
.io_matchBytes_80(matchBytes[80]),
.io_matchBytes_81(matchBytes[81]),
.io_matchBytes_82(matchBytes[82]),
.io_matchBytes_83(matchBytes[83]),
.io_matchBytes_84(matchBytes[84]),
.io_matchBytes_85(matchBytes[85]),
.io_matchBytes_86(matchBytes[86]),
.io_matchBytes_87(matchBytes[87]),
.io_matchBytes_88(matchBytes[88]),
.io_matchBytes_89(matchBytes[89]),
.io_matchBytes_90(matchBytes[90]),
.io_matchBytes_91(matchBytes[91]),
.io_matchBytes_92(matchBytes[92]),
.io_matchBytes_93(matchBytes[93]),
.io_matchBytes_94(matchBytes[94]),
.io_matchBytes_95(matchBytes[95]),
.io_matchBytes_96(matchBytes[96]),
.io_matchBytes_97(matchBytes[97]),
.io_matchBytes_98(matchBytes[98]),
.io_matchBytes_99(matchBytes[99]),
.io_matchBytes_100(matchBytes[100]),
.io_matchBytes_101(matchBytes[101]),
.io_matchBytes_102(matchBytes[102]),
.io_matchBytes_103(matchBytes[103]),
.io_matchBytes_104(matchBytes[104]),
.io_matchBytes_105(matchBytes[105]),
.io_matchBytes_106(matchBytes[106]),
.io_matchBytes_107(matchBytes[107]),
.io_matchBytes_108(matchBytes[108]),
.io_matchBytes_109(matchBytes[109]),
.io_matchBytes_110(matchBytes[110]),
.io_matchBytes_111(matchBytes[111]),
.io_matchBytes_112(matchBytes[112]),
.io_matchBytes_113(matchBytes[113]),
.io_matchBytes_114(matchBytes[114]),
.io_matchBytes_115(matchBytes[115]),
.io_matchBytes_116(matchBytes[116]),
.io_matchBytes_117(matchBytes[117]),
.io_matchBytes_118(matchBytes[118]),
.io_matchBytes_119(matchBytes[119]),
.io_matchBytes_120(matchBytes[120]),
.io_matchBytes_121(matchBytes[121]),
.io_matchBytes_122(matchBytes[122]),
.io_matchBytes_123(matchBytes[123]),
.io_matchBytes_124(matchBytes[124]),
.io_matchBytes_125(matchBytes[125]),
.io_matchBytes_126(matchBytes[126]),
.io_matchBytes_127(matchBytes[127]),
.io_matchBytes_128(matchBytes[128]),
.io_matchBytes_129(matchBytes[129]),
.io_matchBytes_130(matchBytes[130]),
.io_matchBytes_131(matchBytes[131]),
.io_matchBytes_132(matchBytes[132]),
.io_matchBytes_133(matchBytes[133]),
.io_matchBytes_134(matchBytes[134]),
.io_matchBytes_135(matchBytes[135]),
.io_matchBytes_136(matchBytes[136]),
.io_matchBytes_137(matchBytes[137]),
.io_matchBytes_138(matchBytes[138]),
.io_matchBytes_139(matchBytes[139]),
.io_matchBytes_140(matchBytes[140]),
.io_matchBytes_141(matchBytes[141]),
.io_matchBytes_142(matchBytes[142]),
.io_matchBytes_143(matchBytes[143]),
.io_matchBytes_144(matchBytes[144]),
.io_matchBytes_145(matchBytes[145]),
.io_matchBytes_146(matchBytes[146]),
.io_matchBytes_147(matchBytes[147]),
.io_matchBytes_148(matchBytes[148]),
.io_matchBytes_149(matchBytes[149]),
.io_matchBytes_150(matchBytes[150]),
.io_matchBytes_151(matchBytes[151]),
.io_matchBytes_152(matchBytes[152]),
.io_matchBytes_153(matchBytes[153]),
.io_matchBytes_154(matchBytes[154]),
.io_matchBytes_155(matchBytes[155]),
.io_matchBytes_156(matchBytes[156]),
.io_matchBytes_157(matchBytes[157]),
.io_matchBytes_158(matchBytes[158]),
.io_matchBytes_159(matchBytes[159]),
.io_matchBytes_160(matchBytes[160]),
.io_matchBytes_161(matchBytes[161]),
.io_matchBytes_162(matchBytes[162]),
.io_matchBytes_163(matchBytes[163]),
.io_matchBytes_164(matchBytes[164]),
.io_matchBytes_165(matchBytes[165]),
.io_matchBytes_166(matchBytes[166]),
.io_matchBytes_167(matchBytes[167]),
.io_matchBytes_168(matchBytes[168]),
.io_matchBytes_169(matchBytes[169]),
.io_matchBytes_170(matchBytes[170]),
.io_matchBytes_171(matchBytes[171]),
.io_matchBytes_172(matchBytes[172]),
.io_matchBytes_173(matchBytes[173]),
.io_matchBytes_174(matchBytes[174]),
.io_matchBytes_175(matchBytes[175]),
.io_matchBytes_176(matchBytes[176]),
.io_matchBytes_177(matchBytes[177]),
.io_matchBytes_178(matchBytes[178]),
.io_matchBytes_179(matchBytes[179]),
.io_matchBytes_180(matchBytes[180]),
.io_matchBytes_181(matchBytes[181]),
.io_matchBytes_182(matchBytes[182]),
.io_matchBytes_183(matchBytes[183]),
.io_matchBytes_184(matchBytes[184]),
.io_matchBytes_185(matchBytes[185]),
.io_matchBytes_186(matchBytes[186]),
.io_matchBytes_187(matchBytes[187]),
.io_matchBytes_188(matchBytes[188]),
.io_matchBytes_189(matchBytes[189]),
.io_matchBytes_190(matchBytes[190]),
.io_matchBytes_191(matchBytes[191]),
.io_matchBytes_192(matchBytes[192]),
.io_matchBytes_193(matchBytes[193]),
.io_matchBytes_194(matchBytes[194]),
.io_matchBytes_195(matchBytes[195]),
.io_matchBytes_196(matchBytes[196]),
.io_matchBytes_197(matchBytes[197]),
.io_matchBytes_198(matchBytes[198]),
.io_matchBytes_199(matchBytes[199]),
.io_matchBytes_200(matchBytes[200]),
.io_matchBytes_201(matchBytes[201]),
.io_matchBytes_202(matchBytes[202]),
.io_matchBytes_203(matchBytes[203]),
.io_matchBytes_204(matchBytes[204]),
.io_matchBytes_205(matchBytes[205]),
.io_matchBytes_206(matchBytes[206]),
.io_matchBytes_207(matchBytes[207]),
.io_matchBytes_208(matchBytes[208]),
.io_matchBytes_209(matchBytes[209]),
.io_matchBytes_210(matchBytes[210]),
.io_matchBytes_211(matchBytes[211]),
.io_matchBytes_212(matchBytes[212]),
.io_matchBytes_213(matchBytes[213]),
.io_matchBytes_214(matchBytes[214]),
.io_matchBytes_215(matchBytes[215]),
.io_matchBytes_216(matchBytes[216]),
.io_matchBytes_217(matchBytes[217]),
.io_matchBytes_218(matchBytes[218]),
.io_matchBytes_219(matchBytes[219]),
.io_matchBytes_220(matchBytes[220]),
.io_matchBytes_221(matchBytes[221]),
.io_matchBytes_222(matchBytes[222]),
.io_matchBytes_223(matchBytes[223]),
.io_matchBytes_224(matchBytes[224]),
.io_matchBytes_225(matchBytes[225]),
.io_matchBytes_226(matchBytes[226]),
.io_matchBytes_227(matchBytes[227]),
.io_matchBytes_228(matchBytes[228]),
.io_matchBytes_229(matchBytes[229]),
.io_matchBytes_230(matchBytes[230]),
.io_matchBytes_231(matchBytes[231]),
.io_matchBytes_232(matchBytes[232]),
.io_matchBytes_233(matchBytes[233]),
.io_matchBytes_234(matchBytes[234]),
.io_matchBytes_235(matchBytes[235]),
.io_matchBytes_236(matchBytes[236]),
.io_matchBytes_237(matchBytes[237]),
.io_matchBytes_238(matchBytes[238]),
.io_matchBytes_239(matchBytes[239]),
.io_matchBytes_240(matchBytes[240]),
.io_matchBytes_241(matchBytes[241]),
.io_matchBytes_242(matchBytes[242]),
.io_matchBytes_243(matchBytes[243]),
.io_matchBytes_244(matchBytes[244]),
.io_matchBytes_245(matchBytes[245]),
.io_matchBytes_246(matchBytes[246]),
.io_matchBytes_247(matchBytes[247]),
.io_matchBytes_248(matchBytes[248]),
.io_matchBytes_249(matchBytes[249]),
.io_matchBytes_250(matchBytes[250]),
.io_matchBytes_251(matchBytes[251]),
.io_matchBytes_252(matchBytes[252]),
.io_matchBytes_253(matchBytes[253]),
.io_matchBytes_254(matchBytes[254]),
.io_matchBytes_255(matchBytes[255]),
.io_matchBytes_256(matchBytes[256]),
.io_matchBytes_257(matchBytes[257]),
.io_matchBytes_258(matchBytes[258]),
.io_matchBytes_259(matchBytes[259]),
.io_matchBytes_260(matchBytes[260]),
.io_matchBytes_261(matchBytes[261]),
.io_matchBytes_262(matchBytes[262]),
.io_matchBytes_263(matchBytes[263]),
.io_matchBytes_264(matchBytes[264]),
.io_matchBytes_265(matchBytes[265]),
.io_matchBytes_266(matchBytes[266]),
.io_matchBytes_267(matchBytes[267]),
.io_matchBytes_268(matchBytes[268]),
.io_matchBytes_269(matchBytes[269]),
.io_matchBytes_270(matchBytes[270]),
.io_matchBytes_271(matchBytes[271]),
.io_matchBytes_272(matchBytes[272]),
.io_matchBytes_273(matchBytes[273]),
.io_matchBytes_274(matchBytes[274]),
.io_matchBytes_275(matchBytes[275]),
.io_matchBytes_276(matchBytes[276]),
.io_matchBytes_277(matchBytes[277]),
.io_matchBytes_278(matchBytes[278]),
.io_matchBytes_279(matchBytes[279]),
.io_matchBytes_280(matchBytes[280]),
.io_matchBytes_281(matchBytes[281]),
.io_matchBytes_282(matchBytes[282]),
.io_matchBytes_283(matchBytes[283]),
.io_matchBytes_284(matchBytes[284]),
.io_matchBytes_285(matchBytes[285]),
.io_matchBytes_286(matchBytes[286]),
.io_matchBytes_287(matchBytes[287]),
.io_matchBytes_288(matchBytes[288]),
.io_matchBytes_289(matchBytes[289]),
.io_matchBytes_290(matchBytes[290]),
.io_matchBytes_291(matchBytes[291]),
.io_matchBytes_292(matchBytes[292]),
.io_matchBytes_293(matchBytes[293]),
.io_matchBytes_294(matchBytes[294]),
.io_matchBytes_295(matchBytes[295]),
.io_matchBytes_296(matchBytes[296]),
.io_matchBytes_297(matchBytes[297]),
.io_matchBytes_298(matchBytes[298]),
.io_matchBytes_299(matchBytes[299]),
.io_matchBytes_300(matchBytes[300]),
.io_matchBytes_301(matchBytes[301]),
.io_matchBytes_302(matchBytes[302]),
.io_matchBytes_303(matchBytes[303]),
.io_matchBytes_304(matchBytes[304]),
.io_matchBytes_305(matchBytes[305]),
.io_matchBytes_306(matchBytes[306]),
.io_matchBytes_307(matchBytes[307]),
.io_matchBytes_308(matchBytes[308]),
.io_matchBytes_309(matchBytes[309]),
.io_matchBytes_310(matchBytes[310]),
.io_matchBytes_311(matchBytes[311]),
.io_matchBytes_312(matchBytes[312]),
.io_matchBytes_313(matchBytes[313]),
.io_matchBytes_314(matchBytes[314]),
.io_matchBytes_315(matchBytes[315]),
.io_matchBytes_316(matchBytes[316]),
.io_matchBytes_317(matchBytes[317]),
.io_matchBytes_318(matchBytes[318]),
.io_matchBytes_319(matchBytes[319]),
.io_matchBytes_320(matchBytes[320]),
.io_matchBytes_321(matchBytes[321]),
.io_matchBytes_322(matchBytes[322]),
.io_matchBytes_323(matchBytes[323]),
.io_matchBytes_324(matchBytes[324]),
.io_matchBytes_325(matchBytes[325]),
.io_matchBytes_326(matchBytes[326]),
.io_matchBytes_327(matchBytes[327]),
.io_matchBytes_328(matchBytes[328]),
.io_matchBytes_329(matchBytes[329]),
.io_matchBytes_330(matchBytes[330]),
.io_matchBytes_331(matchBytes[331]),
.io_matchBytes_332(matchBytes[332]),
.io_matchBytes_333(matchBytes[333]),
.io_matchBytes_334(matchBytes[334]),
.io_matchBytes_335(matchBytes[335]),
.io_matchBytes_336(matchBytes[336]),
.io_matchBytes_337(matchBytes[337]),
.io_matchBytes_338(matchBytes[338]),
.io_matchBytes_339(matchBytes[339]),
.io_matchBytes_340(matchBytes[340]),
.io_matchBytes_341(matchBytes[341]),
.io_matchBytes_342(matchBytes[342]),
.io_matchBytes_343(matchBytes[343]),
.io_matchBytes_344(matchBytes[344]),
.io_matchBytes_345(matchBytes[345]),
.io_matchBytes_346(matchBytes[346]),
.io_matchBytes_347(matchBytes[347]),
.io_matchBytes_348(matchBytes[348]),
.io_matchBytes_349(matchBytes[349]),
.io_matchBytes_350(matchBytes[350]),
.io_matchBytes_351(matchBytes[351]),
.io_matchBytes_352(matchBytes[352]),
.io_matchBytes_353(matchBytes[353]),
.io_matchBytes_354(matchBytes[354]),
.io_matchBytes_355(matchBytes[355]),
.io_matchBytes_356(matchBytes[356]),
.io_matchBytes_357(matchBytes[357]),
.io_matchBytes_358(matchBytes[358]),
.io_matchBytes_359(matchBytes[359]),
.io_matchBytes_360(matchBytes[360]),
.io_matchBytes_361(matchBytes[361]),
.io_matchBytes_362(matchBytes[362]),
.io_matchBytes_363(matchBytes[363]),
.io_matchBytes_364(matchBytes[364]),
.io_matchBytes_365(matchBytes[365]),
.io_matchBytes_366(matchBytes[366]),
.io_matchBytes_367(matchBytes[367]),
.io_matchBytes_368(matchBytes[368]),
.io_matchBytes_369(matchBytes[369]),
.io_matchBytes_370(matchBytes[370]),
.io_matchBytes_371(matchBytes[371]),
.io_matchBytes_372(matchBytes[372]),
.io_matchBytes_373(matchBytes[373]),
.io_matchBytes_374(matchBytes[374]),
.io_matchBytes_375(matchBytes[375]),
.io_matchBytes_376(matchBytes[376]),
.io_matchBytes_377(matchBytes[377]),
.io_matchBytes_378(matchBytes[378]),
.io_matchBytes_379(matchBytes[379]),
.io_matchBytes_380(matchBytes[380]),
.io_matchBytes_381(matchBytes[381]),
.io_matchBytes_382(matchBytes[382]),
.io_matchBytes_383(matchBytes[383]),
.io_matchBytes_384(matchBytes[384]),
.io_matchBytes_385(matchBytes[385]),
.io_matchBytes_386(matchBytes[386]),
.io_matchBytes_387(matchBytes[387]),
.io_matchBytes_388(matchBytes[388]),
.io_matchBytes_389(matchBytes[389]),
.io_matchBytes_390(matchBytes[390]),
.io_matchBytes_391(matchBytes[391]),
.io_matchBytes_392(matchBytes[392]),
.io_matchBytes_393(matchBytes[393]),
.io_matchBytes_394(matchBytes[394]),
.io_matchBytes_395(matchBytes[395]),
.io_matchBytes_396(matchBytes[396]),
.io_matchBytes_397(matchBytes[397]),
.io_matchBytes_398(matchBytes[398]),
.io_matchBytes_399(matchBytes[399]),
.io_matchBytes_400(matchBytes[400]),
.io_matchBytes_401(matchBytes[401]),
.io_matchBytes_402(matchBytes[402]),
.io_matchBytes_403(matchBytes[403]),
.io_matchBytes_404(matchBytes[404]),
.io_matchBytes_405(matchBytes[405]),
.io_matchBytes_406(matchBytes[406]),
.io_matchBytes_407(matchBytes[407]),
.io_matchBytes_408(matchBytes[408]),
.io_matchBytes_409(matchBytes[409]),
.io_matchBytes_410(matchBytes[410]),
.io_matchBytes_411(matchBytes[411]),
.io_matchBytes_412(matchBytes[412]),
.io_matchBytes_413(matchBytes[413]),
.io_matchBytes_414(matchBytes[414]),
.io_matchBytes_415(matchBytes[415]),
.io_matchBytes_416(matchBytes[416]),
.io_matchBytes_417(matchBytes[417]),
.io_matchBytes_418(matchBytes[418]),
.io_matchBytes_419(matchBytes[419]),
.io_matchBytes_420(matchBytes[420]),
.io_matchBytes_421(matchBytes[421]),
.io_matchBytes_422(matchBytes[422]),
.io_matchBytes_423(matchBytes[423]),
.io_matchBytes_424(matchBytes[424]),
.io_matchBytes_425(matchBytes[425]),
.io_matchBytes_426(matchBytes[426]),
.io_matchBytes_427(matchBytes[427]),
.io_matchBytes_428(matchBytes[428]),
.io_matchBytes_429(matchBytes[429]),
.io_matchBytes_430(matchBytes[430]),
.io_matchBytes_431(matchBytes[431]),
.io_matchBytes_432(matchBytes[432]),
.io_matchBytes_433(matchBytes[433]),
.io_matchBytes_434(matchBytes[434]),
.io_matchBytes_435(matchBytes[435]),
.io_matchBytes_436(matchBytes[436]),
.io_matchBytes_437(matchBytes[437]),
.io_matchBytes_438(matchBytes[438]),
.io_matchBytes_439(matchBytes[439]),
.io_matchBytes_440(matchBytes[440]),
.io_matchBytes_441(matchBytes[441]),
.io_matchBytes_442(matchBytes[442]),
.io_matchBytes_443(matchBytes[443]),
.io_matchBytes_444(matchBytes[444]),
.io_matchBytes_445(matchBytes[445]),
.io_matchBytes_446(matchBytes[446]),
.io_matchBytes_447(matchBytes[447]),
.io_matchBytes_448(matchBytes[448]),
.io_matchBytes_449(matchBytes[449]),
.io_matchBytes_450(matchBytes[450]),
.io_matchBytes_451(matchBytes[451]),
.io_matchBytes_452(matchBytes[452]),
.io_matchBytes_453(matchBytes[453]),
.io_matchBytes_454(matchBytes[454]),
.io_matchBytes_455(matchBytes[455]),
.io_matchBytes_456(matchBytes[456]),
.io_matchBytes_457(matchBytes[457]),
.io_matchBytes_458(matchBytes[458]),
.io_matchBytes_459(matchBytes[459]),
.io_matchBytes_460(matchBytes[460]),
.io_matchBytes_461(matchBytes[461]),
.io_matchBytes_462(matchBytes[462]),
.io_matchBytes_463(matchBytes[463]),
.io_matchBytes_464(matchBytes[464]),
.io_matchBytes_465(matchBytes[465]),
.io_matchBytes_466(matchBytes[466]),
.io_matchBytes_467(matchBytes[467]),
.io_matchBytes_468(matchBytes[468]),
.io_matchBytes_469(matchBytes[469]),
.io_matchBytes_470(matchBytes[470]),
.io_matchBytes_471(matchBytes[471]),
.io_matchBytes_472(matchBytes[472]),
.io_matchBytes_473(matchBytes[473]),
.io_matchBytes_474(matchBytes[474]),
.io_matchBytes_475(matchBytes[475]),
.io_matchBytes_476(matchBytes[476]),
.io_matchBytes_477(matchBytes[477]),
.io_matchBytes_478(matchBytes[478]),
.io_matchBytes_479(matchBytes[479]),
.io_matchBytes_480(matchBytes[480]),
.io_matchBytes_481(matchBytes[481]),
.io_matchBytes_482(matchBytes[482]),
.io_matchBytes_483(matchBytes[483]),
.io_matchBytes_484(matchBytes[484]),
.io_matchBytes_485(matchBytes[485]),
.io_matchBytes_486(matchBytes[486]),
.io_matchBytes_487(matchBytes[487]),
.io_matchBytes_488(matchBytes[488]),
.io_matchBytes_489(matchBytes[489]),
.io_matchBytes_490(matchBytes[490]),
.io_matchBytes_491(matchBytes[491]),
.io_matchBytes_492(matchBytes[492]),
.io_matchBytes_493(matchBytes[493]),
.io_matchBytes_494(matchBytes[494]),
.io_matchBytes_495(matchBytes[495]),
.io_matchBytes_496(matchBytes[496]),
.io_matchBytes_497(matchBytes[497]),
.io_matchBytes_498(matchBytes[498]),
.io_matchBytes_499(matchBytes[499]),
.io_matchBytes_500(matchBytes[500]),
.io_matchBytes_501(matchBytes[501]),
.io_matchBytes_502(matchBytes[502]),
.io_matchBytes_503(matchBytes[503]),
.io_matchBytes_504(matchBytes[504]),
.io_matchBytes_505(matchBytes[505]),
.io_matchBytes_506(matchBytes[506]),
.io_matchBytes_507(matchBytes[507]),
.io_matchBytes_508(matchBytes[508]),
.io_matchBytes_509(matchBytes[509]),
.io_matchBytes_510(matchBytes[510]),
.io_matchBytes_511(matchBytes[511]),
.io_matchBytes_512(matchBytes[512]),
.io_matchBytes_513(matchBytes[513]),
.io_matchBytes_514(matchBytes[514]),
.io_matchBytes_515(matchBytes[515]),
.io_matchBytes_516(matchBytes[516]),
.io_matchBytes_517(matchBytes[517]),
.io_matchBytes_518(matchBytes[518]),
.io_matchBytes_519(matchBytes[519]),
.io_matchBytes_520(matchBytes[520]),
.io_matchBytes_521(matchBytes[521]),
.io_matchBytes_522(matchBytes[522]),
.io_matchBytes_523(matchBytes[523]),
.io_matchBytes_524(matchBytes[524]),
.io_matchBytes_525(matchBytes[525]),
.io_matchBytes_526(matchBytes[526]),
.io_matchBytes_527(matchBytes[527]),
.io_matchBytes_528(matchBytes[528]),
.io_matchBytes_529(matchBytes[529]),
.io_matchBytes_530(matchBytes[530]),
.io_matchBytes_531(matchBytes[531]),
.io_matchBytes_532(matchBytes[532]),
.io_matchBytes_533(matchBytes[533]),
.io_matchBytes_534(matchBytes[534]),
.io_matchBytes_535(matchBytes[535]),
.io_matchBytes_536(matchBytes[536]),
.io_matchBytes_537(matchBytes[537]),
.io_matchBytes_538(matchBytes[538]),
.io_matchBytes_539(matchBytes[539]),
.io_matchBytes_540(matchBytes[540]),
.io_matchBytes_541(matchBytes[541]),
.io_matchBytes_542(matchBytes[542]),
.io_matchBytes_543(matchBytes[543]),
.io_matchBytes_544(matchBytes[544]),
.io_matchBytes_545(matchBytes[545]),
.io_matchBytes_546(matchBytes[546]),
.io_matchBytes_547(matchBytes[547]),
.io_matchBytes_548(matchBytes[548]),
.io_matchBytes_549(matchBytes[549]),
.io_matchBytes_550(matchBytes[550]),
.io_matchBytes_551(matchBytes[551]),
.io_matchBytes_552(matchBytes[552]),
.io_matchBytes_553(matchBytes[553]),
.io_matchBytes_554(matchBytes[554]),
.io_matchBytes_555(matchBytes[555]),
.io_matchBytes_556(matchBytes[556]),
.io_matchBytes_557(matchBytes[557]),
.io_matchBytes_558(matchBytes[558]),
.io_matchBytes_559(matchBytes[559]),
.io_matchBytes_560(matchBytes[560]),
.io_matchBytes_561(matchBytes[561]),
.io_matchBytes_562(matchBytes[562]),
.io_matchBytes_563(matchBytes[563]),
.io_matchBytes_564(matchBytes[564]),
.io_matchBytes_565(matchBytes[565]),
.io_matchBytes_566(matchBytes[566]),
.io_matchBytes_567(matchBytes[567]),
.io_matchBytes_568(matchBytes[568]),
.io_matchBytes_569(matchBytes[569]),
.io_matchBytes_570(matchBytes[570]),
.io_matchBytes_571(matchBytes[571]),
.io_matchBytes_572(matchBytes[572]),
.io_matchBytes_573(matchBytes[573]),
.io_matchBytes_574(matchBytes[574]),
.io_matchBytes_575(matchBytes[575]),
.io_matchBytes_576(matchBytes[576]),
.io_matchBytes_577(matchBytes[577]),
.io_matchBytes_578(matchBytes[578]),
.io_matchBytes_579(matchBytes[579]),
.io_matchBytes_580(matchBytes[580]),
.io_matchBytes_581(matchBytes[581]),
.io_matchBytes_582(matchBytes[582]),
.io_matchBytes_583(matchBytes[583]),
.io_matchBytes_584(matchBytes[584]),
.io_matchBytes_585(matchBytes[585]),
.io_matchBytes_586(matchBytes[586]),
.io_matchBytes_587(matchBytes[587]),
.io_matchBytes_588(matchBytes[588]),
.io_matchBytes_589(matchBytes[589]),
.io_matchBytes_590(matchBytes[590]),
.io_matchBytes_591(matchBytes[591]),
.io_matchBytes_592(matchBytes[592]),
.io_matchBytes_593(matchBytes[593]),
.io_matchBytes_594(matchBytes[594]),
.io_matchBytes_595(matchBytes[595]),
.io_matchBytes_596(matchBytes[596]),
.io_matchBytes_597(matchBytes[597]),
.io_matchBytes_598(matchBytes[598]),
.io_matchBytes_599(matchBytes[599]),
.io_matchBytes_600(matchBytes[600]),
.io_matchBytes_601(matchBytes[601]),
.io_matchBytes_602(matchBytes[602]),
.io_matchBytes_603(matchBytes[603]),
.io_matchBytes_604(matchBytes[604]),
.io_matchBytes_605(matchBytes[605]),
.io_matchBytes_606(matchBytes[606]),
.io_matchBytes_607(matchBytes[607]),
.io_matchBytes_608(matchBytes[608]),
.io_matchBytes_609(matchBytes[609]),
.io_matchBytes_610(matchBytes[610]),
.io_matchBytes_611(matchBytes[611]),
.io_matchBytes_612(matchBytes[612]),
.io_matchBytes_613(matchBytes[613]),
.io_matchBytes_614(matchBytes[614]),
.io_matchBytes_615(matchBytes[615]),
.io_matchBytes_616(matchBytes[616]),
.io_matchBytes_617(matchBytes[617]),
.io_matchBytes_618(matchBytes[618]),
.io_matchBytes_619(matchBytes[619]),
.io_matchBytes_620(matchBytes[620]),
.io_matchBytes_621(matchBytes[621]),
.io_matchBytes_622(matchBytes[622]),
.io_matchBytes_623(matchBytes[623]),
.io_matchBytes_624(matchBytes[624]),
.io_matchBytes_625(matchBytes[625]),
.io_matchBytes_626(matchBytes[626]),
.io_matchBytes_627(matchBytes[627]),
.io_matchBytes_628(matchBytes[628]),
.io_matchBytes_629(matchBytes[629]),
.io_matchBytes_630(matchBytes[630]),
.io_matchBytes_631(matchBytes[631]),
.io_matchBytes_632(matchBytes[632]),
.io_matchBytes_633(matchBytes[633]),
.io_matchBytes_634(matchBytes[634]),
.io_matchBytes_635(matchBytes[635]),
.io_matchBytes_636(matchBytes[636]),
.io_matchBytes_637(matchBytes[637]),
.io_matchBytes_638(matchBytes[638]),
.io_matchBytes_639(matchBytes[639]),
.io_matchBytes_640(matchBytes[640]),
.io_matchBytes_641(matchBytes[641]),
.io_matchBytes_642(matchBytes[642]),
.io_matchBytes_643(matchBytes[643]),
.io_matchBytes_644(matchBytes[644]),
.io_matchBytes_645(matchBytes[645]),
.io_matchBytes_646(matchBytes[646]),
.io_matchBytes_647(matchBytes[647]),
.io_matchBytes_648(matchBytes[648]),
.io_matchBytes_649(matchBytes[649]),
.io_matchBytes_650(matchBytes[650]),
.io_matchBytes_651(matchBytes[651]),
.io_matchBytes_652(matchBytes[652]),
.io_matchBytes_653(matchBytes[653]),
.io_matchBytes_654(matchBytes[654]),
.io_matchBytes_655(matchBytes[655]),
.io_matchBytes_656(matchBytes[656]),
.io_matchBytes_657(matchBytes[657]),
.io_matchBytes_658(matchBytes[658]),
.io_matchBytes_659(matchBytes[659]),
.io_matchBytes_660(matchBytes[660]),
.io_matchBytes_661(matchBytes[661]),
.io_matchBytes_662(matchBytes[662]),
.io_matchBytes_663(matchBytes[663]),
.io_matchBytes_664(matchBytes[664]),
.io_matchBytes_665(matchBytes[665]),
.io_matchBytes_666(matchBytes[666]),
.io_matchBytes_667(matchBytes[667]),
.io_matchBytes_668(matchBytes[668]),
.io_matchBytes_669(matchBytes[669]),
.io_matchBytes_670(matchBytes[670]),
.io_matchBytes_671(matchBytes[671]),
.io_matchBytes_672(matchBytes[672]),
.io_matchBytes_673(matchBytes[673]),
.io_matchBytes_674(matchBytes[674]),
.io_matchBytes_675(matchBytes[675]),
.io_matchBytes_676(matchBytes[676]),
.io_matchBytes_677(matchBytes[677]),
.io_matchBytes_678(matchBytes[678]),
.io_matchBytes_679(matchBytes[679]),
.io_matchBytes_680(matchBytes[680]),
.io_matchBytes_681(matchBytes[681]),
.io_matchBytes_682(matchBytes[682]),
.io_matchBytes_683(matchBytes[683]),
.io_matchBytes_684(matchBytes[684]),
.io_matchBytes_685(matchBytes[685]),
.io_matchBytes_686(matchBytes[686]),
.io_matchBytes_687(matchBytes[687]),
.io_matchBytes_688(matchBytes[688]),
.io_matchBytes_689(matchBytes[689]),
.io_matchBytes_690(matchBytes[690]),
.io_matchBytes_691(matchBytes[691]),
.io_matchBytes_692(matchBytes[692]),
.io_matchBytes_693(matchBytes[693]),
.io_matchBytes_694(matchBytes[694]),
.io_matchBytes_695(matchBytes[695]),
.io_matchBytes_696(matchBytes[696]),
.io_matchBytes_697(matchBytes[697]),
.io_matchBytes_698(matchBytes[698]),
.io_matchBytes_699(matchBytes[699]),
.io_matchBytes_700(matchBytes[700]),
.io_matchBytes_701(matchBytes[701]),
.io_matchBytes_702(matchBytes[702]),
.io_matchBytes_703(matchBytes[703]),
.io_matchBytes_704(matchBytes[704]),
.io_matchBytes_705(matchBytes[705]),
.io_matchBytes_706(matchBytes[706]),
.io_matchBytes_707(matchBytes[707]),
.io_matchBytes_708(matchBytes[708]),
.io_matchBytes_709(matchBytes[709]),
.io_matchBytes_710(matchBytes[710]),
.io_matchBytes_711(matchBytes[711]),
.io_matchBytes_712(matchBytes[712]),
.io_matchBytes_713(matchBytes[713]),
.io_matchBytes_714(matchBytes[714]),
.io_matchBytes_715(matchBytes[715]),
.io_matchBytes_716(matchBytes[716]),
.io_matchBytes_717(matchBytes[717]),
.io_matchBytes_718(matchBytes[718]),
.io_matchBytes_719(matchBytes[719]),
.io_matchBytes_720(matchBytes[720]),
.io_matchBytes_721(matchBytes[721]),
.io_matchBytes_722(matchBytes[722]),
.io_matchBytes_723(matchBytes[723]),
.io_matchBytes_724(matchBytes[724]),
.io_matchBytes_725(matchBytes[725]),
.io_matchBytes_726(matchBytes[726]),
.io_matchBytes_727(matchBytes[727]),
.io_matchBytes_728(matchBytes[728]),
.io_matchBytes_729(matchBytes[729]),
.io_matchBytes_730(matchBytes[730]),
.io_matchBytes_731(matchBytes[731]),
.io_matchBytes_732(matchBytes[732]),
.io_matchBytes_733(matchBytes[733]),
.io_matchBytes_734(matchBytes[734]),
.io_matchBytes_735(matchBytes[735]),
.io_matchBytes_736(matchBytes[736]),
.io_matchBytes_737(matchBytes[737]),
.io_matchBytes_738(matchBytes[738]),
.io_matchBytes_739(matchBytes[739]),
.io_matchBytes_740(matchBytes[740]),
.io_matchBytes_741(matchBytes[741]),
.io_matchBytes_742(matchBytes[742]),
.io_matchBytes_743(matchBytes[743]),
.io_matchBytes_744(matchBytes[744]),
.io_matchBytes_745(matchBytes[745]),
.io_matchBytes_746(matchBytes[746]),
.io_matchBytes_747(matchBytes[747]),
.io_matchBytes_748(matchBytes[748]),
.io_matchBytes_749(matchBytes[749]),
.io_matchBytes_750(matchBytes[750]),
.io_matchBytes_751(matchBytes[751]),
.io_matchBytes_752(matchBytes[752]),
.io_matchBytes_753(matchBytes[753]),
.io_matchBytes_754(matchBytes[754]),
.io_matchBytes_755(matchBytes[755]),
.io_matchBytes_756(matchBytes[756]),
.io_matchBytes_757(matchBytes[757]),
.io_matchBytes_758(matchBytes[758]),
.io_matchBytes_759(matchBytes[759]),
.io_matchBytes_760(matchBytes[760]),
.io_matchBytes_761(matchBytes[761]),
.io_matchBytes_762(matchBytes[762]),
.io_matchBytes_763(matchBytes[763]),
.io_matchBytes_764(matchBytes[764]),
.io_matchBytes_765(matchBytes[765]),
.io_matchBytes_766(matchBytes[766]),
.io_matchBytes_767(matchBytes[767]),
.io_matchBytes_768(matchBytes[768]),
.io_matchBytes_769(matchBytes[769]),
.io_matchBytes_770(matchBytes[770]),
.io_matchBytes_771(matchBytes[771]),
.io_matchBytes_772(matchBytes[772]),
.io_matchBytes_773(matchBytes[773]),
.io_matchBytes_774(matchBytes[774]),
.io_matchBytes_775(matchBytes[775]),
.io_matchBytes_776(matchBytes[776]),
.io_matchBytes_777(matchBytes[777]),
.io_matchBytes_778(matchBytes[778]),
.io_matchBytes_779(matchBytes[779]),
.io_matchBytes_780(matchBytes[780]),
.io_matchBytes_781(matchBytes[781]),
.io_matchBytes_782(matchBytes[782]),
.io_matchBytes_783(matchBytes[783]),
.io_matchBytes_784(matchBytes[784]),
.io_matchBytes_785(matchBytes[785]),
.io_matchBytes_786(matchBytes[786]),
.io_matchBytes_787(matchBytes[787]),
.io_matchBytes_788(matchBytes[788]),
.io_matchBytes_789(matchBytes[789]),
.io_matchBytes_790(matchBytes[790]),
.io_matchBytes_791(matchBytes[791]),
.io_matchBytes_792(matchBytes[792]),
.io_matchBytes_793(matchBytes[793]),
.io_matchBytes_794(matchBytes[794]),
.io_matchBytes_795(matchBytes[795]),
.io_matchBytes_796(matchBytes[796]),
.io_matchBytes_797(matchBytes[797]),
.io_matchBytes_798(matchBytes[798]),
.io_matchBytes_799(matchBytes[799]),
.io_matchBytes_800(matchBytes[800]),
.io_matchBytes_801(matchBytes[801]),
.io_matchBytes_802(matchBytes[802]),
.io_matchBytes_803(matchBytes[803]),
.io_matchBytes_804(matchBytes[804]),
.io_matchBytes_805(matchBytes[805]),
.io_matchBytes_806(matchBytes[806]),
.io_matchBytes_807(matchBytes[807]),
.io_matchBytes_808(matchBytes[808]),
.io_matchBytes_809(matchBytes[809]),
.io_matchBytes_810(matchBytes[810]),
.io_matchBytes_811(matchBytes[811]),
.io_matchBytes_812(matchBytes[812]),
.io_matchBytes_813(matchBytes[813]),
.io_matchBytes_814(matchBytes[814]),
.io_matchBytes_815(matchBytes[815]),
.io_matchBytes_816(matchBytes[816]),
.io_matchBytes_817(matchBytes[817]),
.io_matchBytes_818(matchBytes[818]),
.io_matchBytes_819(matchBytes[819]),
.io_matchBytes_820(matchBytes[820]),
.io_matchBytes_821(matchBytes[821]),
.io_matchBytes_822(matchBytes[822]),
.io_matchBytes_823(matchBytes[823]),
.io_matchBytes_824(matchBytes[824]),
.io_matchBytes_825(matchBytes[825]),
.io_matchBytes_826(matchBytes[826]),
.io_matchBytes_827(matchBytes[827]),
.io_matchBytes_828(matchBytes[828]),
.io_matchBytes_829(matchBytes[829]),
.io_matchBytes_830(matchBytes[830]),
.io_matchBytes_831(matchBytes[831]),
.io_matchBytes_832(matchBytes[832]),
.io_matchBytes_833(matchBytes[833]),
.io_matchBytes_834(matchBytes[834]),
.io_matchBytes_835(matchBytes[835]),
.io_matchBytes_836(matchBytes[836]),
.io_matchBytes_837(matchBytes[837]),
.io_matchBytes_838(matchBytes[838]),
.io_matchBytes_839(matchBytes[839]),
.io_matchBytes_840(matchBytes[840]),
.io_matchBytes_841(matchBytes[841]),
.io_matchBytes_842(matchBytes[842]),
.io_matchBytes_843(matchBytes[843]),
.io_matchBytes_844(matchBytes[844]),
.io_matchBytes_845(matchBytes[845]),
.io_matchBytes_846(matchBytes[846]),
.io_matchBytes_847(matchBytes[847]),
.io_matchBytes_848(matchBytes[848]),
.io_matchBytes_849(matchBytes[849]),
.io_matchBytes_850(matchBytes[850]),
.io_matchBytes_851(matchBytes[851]),
.io_matchBytes_852(matchBytes[852]),
.io_matchBytes_853(matchBytes[853]),
.io_matchBytes_854(matchBytes[854]),
.io_matchBytes_855(matchBytes[855]),
.io_matchBytes_856(matchBytes[856]),
.io_matchBytes_857(matchBytes[857]),
.io_matchBytes_858(matchBytes[858]),
.io_matchBytes_859(matchBytes[859]),
.io_matchBytes_860(matchBytes[860]),
.io_matchBytes_861(matchBytes[861]),
.io_matchBytes_862(matchBytes[862]),
.io_matchBytes_863(matchBytes[863]),
.io_matchBytes_864(matchBytes[864]),
.io_matchBytes_865(matchBytes[865]),
.io_matchBytes_866(matchBytes[866]),
.io_matchBytes_867(matchBytes[867]),
.io_matchBytes_868(matchBytes[868]),
.io_matchBytes_869(matchBytes[869]),
.io_matchBytes_870(matchBytes[870]),
.io_matchBytes_871(matchBytes[871]),
.io_matchBytes_872(matchBytes[872]),
.io_matchBytes_873(matchBytes[873]),
.io_matchBytes_874(matchBytes[874]),
.io_matchBytes_875(matchBytes[875]),
.io_matchBytes_876(matchBytes[876]),
.io_matchBytes_877(matchBytes[877]),
.io_matchBytes_878(matchBytes[878]),
.io_matchBytes_879(matchBytes[879]),
.io_matchBytes_880(matchBytes[880]),
.io_matchBytes_881(matchBytes[881]),
.io_matchBytes_882(matchBytes[882]),
.io_matchBytes_883(matchBytes[883]),
.io_matchBytes_884(matchBytes[884]),
.io_matchBytes_885(matchBytes[885]),
.io_matchBytes_886(matchBytes[886]),
.io_matchBytes_887(matchBytes[887]),
.io_matchBytes_888(matchBytes[888]),
.io_matchBytes_889(matchBytes[889]),
.io_matchBytes_890(matchBytes[890]),
.io_matchBytes_891(matchBytes[891]),
.io_matchBytes_892(matchBytes[892]),
.io_matchBytes_893(matchBytes[893]),
.io_matchBytes_894(matchBytes[894]),
.io_matchBytes_895(matchBytes[895]),
.io_matchBytes_896(matchBytes[896]),
.io_matchBytes_897(matchBytes[897]),
.io_matchBytes_898(matchBytes[898]),
.io_matchBytes_899(matchBytes[899]),
.io_matchBytes_900(matchBytes[900]),
.io_matchBytes_901(matchBytes[901]),
.io_matchBytes_902(matchBytes[902]),
.io_matchBytes_903(matchBytes[903]),
.io_matchBytes_904(matchBytes[904]),
.io_matchBytes_905(matchBytes[905]),
.io_matchBytes_906(matchBytes[906]),
.io_matchBytes_907(matchBytes[907]),
.io_matchBytes_908(matchBytes[908]),
.io_matchBytes_909(matchBytes[909]),
.io_matchBytes_910(matchBytes[910]),
.io_matchBytes_911(matchBytes[911]),
.io_matchBytes_912(matchBytes[912]),
.io_matchBytes_913(matchBytes[913]),
.io_matchBytes_914(matchBytes[914]),
.io_matchBytes_915(matchBytes[915]),
.io_matchBytes_916(matchBytes[916]),
.io_matchBytes_917(matchBytes[917]),
.io_matchBytes_918(matchBytes[918]),
.io_matchBytes_919(matchBytes[919]),
.io_matchBytes_920(matchBytes[920]),
.io_matchBytes_921(matchBytes[921]),
.io_matchBytes_922(matchBytes[922]),
.io_matchBytes_923(matchBytes[923]),
.io_matchBytes_924(matchBytes[924]),
.io_matchBytes_925(matchBytes[925]),
.io_matchBytes_926(matchBytes[926]),
.io_matchBytes_927(matchBytes[927]),
.io_matchBytes_928(matchBytes[928]),
.io_matchBytes_929(matchBytes[929]),
.io_matchBytes_930(matchBytes[930]),
.io_matchBytes_931(matchBytes[931]),
.io_matchBytes_932(matchBytes[932]),
.io_matchBytes_933(matchBytes[933]),
.io_matchBytes_934(matchBytes[934]),
.io_matchBytes_935(matchBytes[935]),
.io_matchBytes_936(matchBytes[936]),
.io_matchBytes_937(matchBytes[937]),
.io_matchBytes_938(matchBytes[938]),
.io_matchBytes_939(matchBytes[939]),
.io_matchBytes_940(matchBytes[940]),
.io_matchBytes_941(matchBytes[941]),
.io_matchBytes_942(matchBytes[942]),
.io_matchBytes_943(matchBytes[943]),
.io_matchBytes_944(matchBytes[944]),
.io_matchBytes_945(matchBytes[945]),
.io_matchBytes_946(matchBytes[946]),
.io_matchBytes_947(matchBytes[947]),
.io_matchBytes_948(matchBytes[948]),
.io_matchBytes_949(matchBytes[949]),
.io_matchBytes_950(matchBytes[950]),
.io_matchBytes_951(matchBytes[951]),
.io_matchBytes_952(matchBytes[952]),
.io_matchBytes_953(matchBytes[953]),
.io_matchBytes_954(matchBytes[954]),
.io_matchBytes_955(matchBytes[955]),
.io_matchBytes_956(matchBytes[956]),
.io_matchBytes_957(matchBytes[957]),
.io_matchBytes_958(matchBytes[958]),
.io_matchBytes_959(matchBytes[959]),
.io_matchBytes_960(matchBytes[960]),
.io_matchBytes_961(matchBytes[961]),
.io_matchBytes_962(matchBytes[962]),
.io_matchBytes_963(matchBytes[963]),
.io_matchBytes_964(matchBytes[964]),
.io_matchBytes_965(matchBytes[965]),
.io_matchBytes_966(matchBytes[966]),
.io_matchBytes_967(matchBytes[967]),
.io_matchBytes_968(matchBytes[968]),
.io_matchBytes_969(matchBytes[969]),
.io_matchBytes_970(matchBytes[970]),
.io_matchBytes_971(matchBytes[971]),
.io_matchBytes_972(matchBytes[972]),
.io_matchBytes_973(matchBytes[973]),
.io_matchBytes_974(matchBytes[974]),
.io_matchBytes_975(matchBytes[975]),
.io_matchBytes_976(matchBytes[976]),
.io_matchBytes_977(matchBytes[977]),
.io_matchBytes_978(matchBytes[978]),
.io_matchBytes_979(matchBytes[979]),
.io_matchBytes_980(matchBytes[980]),
.io_matchBytes_981(matchBytes[981]),
.io_matchBytes_982(matchBytes[982]),
.io_matchBytes_983(matchBytes[983]),
.io_matchBytes_984(matchBytes[984]),
.io_matchBytes_985(matchBytes[985]),
.io_matchBytes_986(matchBytes[986]),
.io_matchBytes_987(matchBytes[987]),
.io_matchBytes_988(matchBytes[988]),
.io_matchBytes_989(matchBytes[989]),
.io_matchBytes_990(matchBytes[990]),
.io_matchBytes_991(matchBytes[991]),
.io_matchBytes_992(matchBytes[992]),
.io_matchBytes_993(matchBytes[993]),
.io_matchBytes_994(matchBytes[994]),
.io_matchBytes_995(matchBytes[995]),
.io_matchBytes_996(matchBytes[996]),
.io_matchBytes_997(matchBytes[997]),
.io_matchBytes_998(matchBytes[998]),
.io_matchBytes_999(matchBytes[999]),
.io_matchBytes_1000(matchBytes[1000]),
.io_matchBytes_1001(matchBytes[1001]),
.io_matchBytes_1002(matchBytes[1002]),
.io_matchBytes_1003(matchBytes[1003]),
.io_matchBytes_1004(matchBytes[1004]),
.io_matchBytes_1005(matchBytes[1005]),
.io_matchBytes_1006(matchBytes[1006]),
.io_matchBytes_1007(matchBytes[1007]),
.io_matchBytes_1008(matchBytes[1008]),
.io_matchBytes_1009(matchBytes[1009]),
.io_matchBytes_1010(matchBytes[1010]),
.io_matchBytes_1011(matchBytes[1011]),
.io_matchBytes_1012(matchBytes[1012]),
.io_matchBytes_1013(matchBytes[1013]),
.io_matchBytes_1014(matchBytes[1014]),
.io_matchBytes_1015(matchBytes[1015]),
.io_matchBytes_1016(matchBytes[1016]),
.io_matchBytes_1017(matchBytes[1017]),
.io_matchBytes_1018(matchBytes[1018]),
.io_matchBytes_1019(matchBytes[1019]),
.io_matchBytes_1020(matchBytes[1020]),
.io_matchBytes_1021(matchBytes[1021]),
.io_matchBytes_1022(matchBytes[1022]),
.io_matchBytes_1023(matchBytes[1023]),
.io_matchBytes_1024(matchBytes[1024]),
.io_matchBytes_1025(matchBytes[1025]),
.io_matchBytes_1026(matchBytes[1026]),
.io_matchBytes_1027(matchBytes[1027]),
.io_matchBytes_1028(matchBytes[1028]),
.io_matchBytes_1029(matchBytes[1029]),
.io_matchBytes_1030(matchBytes[1030]),
.io_matchBytes_1031(matchBytes[1031]),
.io_matchBytes_1032(matchBytes[1032]),
.io_matchBytes_1033(matchBytes[1033]),
.io_matchBytes_1034(matchBytes[1034]),
.io_matchBytes_1035(matchBytes[1035]),
.io_matchBytes_1036(matchBytes[1036]),
.io_matchBytes_1037(matchBytes[1037]),
.io_matchBytes_1038(matchBytes[1038]),
.io_matchBytes_1039(matchBytes[1039]),
.io_matchBytes_1040(matchBytes[1040]),
.io_matchBytes_1041(matchBytes[1041]),
.io_matchBytes_1042(matchBytes[1042]),
.io_matchBytes_1043(matchBytes[1043]),
.io_matchBytes_1044(matchBytes[1044]),
.io_matchBytes_1045(matchBytes[1045]),
.io_matchBytes_1046(matchBytes[1046]),
.io_matchBytes_1047(matchBytes[1047]),
.io_matchBytes_1048(matchBytes[1048]),
.io_matchBytes_1049(matchBytes[1049]),
.io_matchBytes_1050(matchBytes[1050]),
.io_matchBytes_1051(matchBytes[1051]),
.io_matchBytes_1052(matchBytes[1052]),
.io_matchBytes_1053(matchBytes[1053]),
.io_matchBytes_1054(matchBytes[1054]),
.io_matchBytes_1055(matchBytes[1055]),
.io_matchBytes_1056(matchBytes[1056]),
.io_matchBytes_1057(matchBytes[1057]),
.io_matchBytes_1058(matchBytes[1058]),
.io_matchBytes_1059(matchBytes[1059]),
.io_matchBytes_1060(matchBytes[1060]),
.io_matchBytes_1061(matchBytes[1061]),
.io_matchBytes_1062(matchBytes[1062]),
.io_matchBytes_1063(matchBytes[1063]),
.io_matchBytes_1064(matchBytes[1064]),
.io_matchBytes_1065(matchBytes[1065]),
.io_matchBytes_1066(matchBytes[1066]),
.io_matchBytes_1067(matchBytes[1067]),
.io_matchBytes_1068(matchBytes[1068]),
.io_matchBytes_1069(matchBytes[1069]),
.io_matchBytes_1070(matchBytes[1070]),
.io_matchBytes_1071(matchBytes[1071]),
.io_matchBytes_1072(matchBytes[1072]),
.io_matchBytes_1073(matchBytes[1073]),
.io_matchBytes_1074(matchBytes[1074]),
.io_matchBytes_1075(matchBytes[1075]),
.io_matchBytes_1076(matchBytes[1076]),
.io_matchBytes_1077(matchBytes[1077]),
.io_matchBytes_1078(matchBytes[1078]),
.io_matchBytes_1079(matchBytes[1079]),
.io_matchBytes_1080(matchBytes[1080]),
.io_matchBytes_1081(matchBytes[1081]),
.io_matchBytes_1082(matchBytes[1082]),
.io_matchBytes_1083(matchBytes[1083]),
.io_matchBytes_1084(matchBytes[1084]),
.io_matchBytes_1085(matchBytes[1085]),
.io_matchBytes_1086(matchBytes[1086]),
.io_matchBytes_1087(matchBytes[1087]),
.io_matchBytes_1088(matchBytes[1088]),
.io_matchBytes_1089(matchBytes[1089]),
.io_matchBytes_1090(matchBytes[1090]),
.io_matchBytes_1091(matchBytes[1091]),
.io_matchBytes_1092(matchBytes[1092]),
.io_matchBytes_1093(matchBytes[1093]),
.io_matchBytes_1094(matchBytes[1094]),
.io_matchBytes_1095(matchBytes[1095]),
.io_matchBytes_1096(matchBytes[1096]),
.io_matchBytes_1097(matchBytes[1097]),
.io_matchBytes_1098(matchBytes[1098]),
.io_matchBytes_1099(matchBytes[1099]),
.io_matchBytes_1100(matchBytes[1100]),
.io_matchBytes_1101(matchBytes[1101]),
.io_matchBytes_1102(matchBytes[1102]),
.io_matchBytes_1103(matchBytes[1103]),
.io_matchBytes_1104(matchBytes[1104]),
.io_matchBytes_1105(matchBytes[1105]),
.io_matchBytes_1106(matchBytes[1106]),
.io_matchBytes_1107(matchBytes[1107]),
.io_matchBytes_1108(matchBytes[1108]),
.io_matchBytes_1109(matchBytes[1109]),
.io_matchBytes_1110(matchBytes[1110]),
.io_matchBytes_1111(matchBytes[1111]),
.io_matchBytes_1112(matchBytes[1112]),
.io_matchBytes_1113(matchBytes[1113]),
.io_matchBytes_1114(matchBytes[1114]),
.io_matchBytes_1115(matchBytes[1115]),
.io_matchBytes_1116(matchBytes[1116]),
.io_matchBytes_1117(matchBytes[1117]),
.io_matchBytes_1118(matchBytes[1118]),
.io_matchBytes_1119(matchBytes[1119]),
.io_matchBytes_1120(matchBytes[1120]),
.io_matchBytes_1121(matchBytes[1121]),
.io_matchBytes_1122(matchBytes[1122]),
.io_matchBytes_1123(matchBytes[1123]),
.io_matchBytes_1124(matchBytes[1124]),
.io_matchBytes_1125(matchBytes[1125]),
.io_matchBytes_1126(matchBytes[1126]),
.io_matchBytes_1127(matchBytes[1127]),
.io_matchBytes_1128(matchBytes[1128]),
.io_matchBytes_1129(matchBytes[1129]),
.io_matchBytes_1130(matchBytes[1130]),
.io_matchBytes_1131(matchBytes[1131]),
.io_matchBytes_1132(matchBytes[1132]),
.io_matchBytes_1133(matchBytes[1133]),
.io_matchBytes_1134(matchBytes[1134]),
.io_matchBytes_1135(matchBytes[1135]),
.io_matchBytes_1136(matchBytes[1136]),
.io_matchBytes_1137(matchBytes[1137]),
.io_matchBytes_1138(matchBytes[1138]),
.io_matchBytes_1139(matchBytes[1139]),
.io_matchBytes_1140(matchBytes[1140]),
.io_matchBytes_1141(matchBytes[1141]),
.io_matchBytes_1142(matchBytes[1142]),
.io_matchBytes_1143(matchBytes[1143]),
.io_matchBytes_1144(matchBytes[1144]),
.io_matchBytes_1145(matchBytes[1145]),
.io_matchBytes_1146(matchBytes[1146]),
.io_matchBytes_1147(matchBytes[1147]),
.io_matchBytes_1148(matchBytes[1148]),
.io_matchBytes_1149(matchBytes[1149]),
.io_matchBytes_1150(matchBytes[1150]),
.io_matchBytes_1151(matchBytes[1151]),
.io_matchBytes_1152(matchBytes[1152]),
.io_matchBytes_1153(matchBytes[1153]),
.io_matchBytes_1154(matchBytes[1154]),
.io_matchBytes_1155(matchBytes[1155]),
.io_matchBytes_1156(matchBytes[1156]),
.io_matchBytes_1157(matchBytes[1157]),
.io_matchBytes_1158(matchBytes[1158]),
.io_matchBytes_1159(matchBytes[1159]),
.io_matchBytes_1160(matchBytes[1160]),
.io_matchBytes_1161(matchBytes[1161]),
.io_matchBytes_1162(matchBytes[1162]),
.io_matchBytes_1163(matchBytes[1163]),
.io_matchBytes_1164(matchBytes[1164]),
.io_matchBytes_1165(matchBytes[1165]),
.io_matchBytes_1166(matchBytes[1166]),
.io_matchBytes_1167(matchBytes[1167]),
.io_matchBytes_1168(matchBytes[1168]),
.io_matchBytes_1169(matchBytes[1169]),
.io_matchBytes_1170(matchBytes[1170]),
.io_matchBytes_1171(matchBytes[1171]),
.io_matchBytes_1172(matchBytes[1172]),
.io_matchBytes_1173(matchBytes[1173]),
.io_matchBytes_1174(matchBytes[1174]),
.io_matchBytes_1175(matchBytes[1175]),
.io_matchBytes_1176(matchBytes[1176]),
.io_matchBytes_1177(matchBytes[1177]),
.io_matchBytes_1178(matchBytes[1178]),
.io_matchBytes_1179(matchBytes[1179]),
.io_matchBytes_1180(matchBytes[1180]),
.io_matchBytes_1181(matchBytes[1181]),
.io_matchBytes_1182(matchBytes[1182]),
.io_matchBytes_1183(matchBytes[1183]),
.io_matchBytes_1184(matchBytes[1184]),
.io_matchBytes_1185(matchBytes[1185]),
.io_matchBytes_1186(matchBytes[1186]),
.io_matchBytes_1187(matchBytes[1187]),
.io_matchBytes_1188(matchBytes[1188]),
.io_matchBytes_1189(matchBytes[1189]),
.io_matchBytes_1190(matchBytes[1190]),
.io_matchBytes_1191(matchBytes[1191]),
.io_matchBytes_1192(matchBytes[1192]),
.io_matchBytes_1193(matchBytes[1193]),
.io_matchBytes_1194(matchBytes[1194]),
.io_matchBytes_1195(matchBytes[1195]),
.io_matchBytes_1196(matchBytes[1196]),
.io_matchBytes_1197(matchBytes[1197]),
.io_matchBytes_1198(matchBytes[1198]),
.io_matchBytes_1199(matchBytes[1199]),
.io_matchBytes_1200(matchBytes[1200]),
.io_matchBytes_1201(matchBytes[1201]),
.io_matchBytes_1202(matchBytes[1202]),
.io_matchBytes_1203(matchBytes[1203]),
.io_matchBytes_1204(matchBytes[1204]),
.io_matchBytes_1205(matchBytes[1205]),
.io_matchBytes_1206(matchBytes[1206]),
.io_matchBytes_1207(matchBytes[1207]),
.io_matchBytes_1208(matchBytes[1208]),
.io_matchBytes_1209(matchBytes[1209]),
.io_matchBytes_1210(matchBytes[1210]),
.io_matchBytes_1211(matchBytes[1211]),
.io_matchBytes_1212(matchBytes[1212]),
.io_matchBytes_1213(matchBytes[1213]),
.io_matchBytes_1214(matchBytes[1214]),
.io_matchBytes_1215(matchBytes[1215]),
.io_matchBytes_1216(matchBytes[1216]),
.io_matchBytes_1217(matchBytes[1217]),
.io_matchBytes_1218(matchBytes[1218]),
.io_matchBytes_1219(matchBytes[1219]),
.io_matchBytes_1220(matchBytes[1220]),
.io_matchBytes_1221(matchBytes[1221]),
.io_matchBytes_1222(matchBytes[1222]),
.io_matchBytes_1223(matchBytes[1223]),
.io_matchBytes_1224(matchBytes[1224]),
.io_matchBytes_1225(matchBytes[1225]),
.io_matchBytes_1226(matchBytes[1226]),
.io_matchBytes_1227(matchBytes[1227]),
.io_matchBytes_1228(matchBytes[1228]),
.io_matchBytes_1229(matchBytes[1229]),
.io_matchBytes_1230(matchBytes[1230]),
.io_matchBytes_1231(matchBytes[1231]),
.io_matchBytes_1232(matchBytes[1232]),
.io_matchBytes_1233(matchBytes[1233]),
.io_matchBytes_1234(matchBytes[1234]),
.io_matchBytes_1235(matchBytes[1235]),
.io_matchBytes_1236(matchBytes[1236]),
.io_matchBytes_1237(matchBytes[1237]),
.io_matchBytes_1238(matchBytes[1238]),
.io_matchBytes_1239(matchBytes[1239]),
.io_matchBytes_1240(matchBytes[1240]),
.io_matchBytes_1241(matchBytes[1241]),
.io_matchBytes_1242(matchBytes[1242]),
.io_matchBytes_1243(matchBytes[1243]),
.io_matchBytes_1244(matchBytes[1244]),
.io_matchBytes_1245(matchBytes[1245]),
.io_matchBytes_1246(matchBytes[1246]),
.io_matchBytes_1247(matchBytes[1247]),
.io_matchBytes_1248(matchBytes[1248]),
.io_matchBytes_1249(matchBytes[1249]),
.io_matchBytes_1250(matchBytes[1250]),
.io_matchBytes_1251(matchBytes[1251]),
.io_matchBytes_1252(matchBytes[1252]),
.io_matchBytes_1253(matchBytes[1253]),
.io_matchBytes_1254(matchBytes[1254]),
.io_matchBytes_1255(matchBytes[1255]),
.io_matchBytes_1256(matchBytes[1256]),
.io_matchBytes_1257(matchBytes[1257]),
.io_matchBytes_1258(matchBytes[1258]),
.io_matchBytes_1259(matchBytes[1259]),
.io_matchBytes_1260(matchBytes[1260]),
.io_matchBytes_1261(matchBytes[1261]),
.io_matchBytes_1262(matchBytes[1262]),
.io_matchBytes_1263(matchBytes[1263]),
.io_matchBytes_1264(matchBytes[1264]),
.io_matchBytes_1265(matchBytes[1265]),
.io_matchBytes_1266(matchBytes[1266]),
.io_matchBytes_1267(matchBytes[1267]),
.io_matchBytes_1268(matchBytes[1268]),
.io_matchBytes_1269(matchBytes[1269]),
.io_matchBytes_1270(matchBytes[1270]),
.io_matchBytes_1271(matchBytes[1271]),
.io_matchBytes_1272(matchBytes[1272]),
.io_matchBytes_1273(matchBytes[1273]),
.io_matchBytes_1274(matchBytes[1274]),
.io_matchBytes_1275(matchBytes[1275]),
.io_matchBytes_1276(matchBytes[1276]),
.io_matchBytes_1277(matchBytes[1277]),
.io_matchBytes_1278(matchBytes[1278]),
.io_matchBytes_1279(matchBytes[1279]),
.io_matchBytes_1280(matchBytes[1280]),
.io_matchBytes_1281(matchBytes[1281]),
.io_matchBytes_1282(matchBytes[1282]),
.io_matchBytes_1283(matchBytes[1283]),
.io_matchBytes_1284(matchBytes[1284]),
.io_matchBytes_1285(matchBytes[1285]),
.io_matchBytes_1286(matchBytes[1286]),
.io_matchBytes_1287(matchBytes[1287]),
.io_matchBytes_1288(matchBytes[1288]),
.io_matchBytes_1289(matchBytes[1289]),
.io_matchBytes_1290(matchBytes[1290]),
.io_matchBytes_1291(matchBytes[1291]),
.io_matchBytes_1292(matchBytes[1292]),
.io_matchBytes_1293(matchBytes[1293]),
.io_matchBytes_1294(matchBytes[1294]),
.io_matchBytes_1295(matchBytes[1295]),
.io_matchBytes_1296(matchBytes[1296]),
.io_matchBytes_1297(matchBytes[1297]),
.io_matchBytes_1298(matchBytes[1298]),
.io_matchBytes_1299(matchBytes[1299]),
.io_matchBytes_1300(matchBytes[1300]),
.io_matchBytes_1301(matchBytes[1301]),
.io_matchBytes_1302(matchBytes[1302]),
.io_matchBytes_1303(matchBytes[1303]),
.io_matchBytes_1304(matchBytes[1304]),
.io_matchBytes_1305(matchBytes[1305]),
.io_matchBytes_1306(matchBytes[1306]),
.io_matchBytes_1307(matchBytes[1307]),
.io_matchBytes_1308(matchBytes[1308]),
.io_matchBytes_1309(matchBytes[1309]),
.io_matchBytes_1310(matchBytes[1310]),
.io_matchBytes_1311(matchBytes[1311]),
.io_matchBytes_1312(matchBytes[1312]),
.io_matchBytes_1313(matchBytes[1313]),
.io_matchBytes_1314(matchBytes[1314]),
.io_matchBytes_1315(matchBytes[1315]),
.io_matchBytes_1316(matchBytes[1316]),
.io_matchBytes_1317(matchBytes[1317]),
.io_matchBytes_1318(matchBytes[1318]),
.io_matchBytes_1319(matchBytes[1319]),
.io_matchBytes_1320(matchBytes[1320]),
.io_matchBytes_1321(matchBytes[1321]),
.io_matchBytes_1322(matchBytes[1322]),
.io_matchBytes_1323(matchBytes[1323]),
.io_matchBytes_1324(matchBytes[1324]),
.io_matchBytes_1325(matchBytes[1325]),
.io_matchBytes_1326(matchBytes[1326]),
.io_matchBytes_1327(matchBytes[1327]),
.io_matchBytes_1328(matchBytes[1328]),
.io_matchBytes_1329(matchBytes[1329]),
.io_matchBytes_1330(matchBytes[1330]),
.io_matchBytes_1331(matchBytes[1331]),
.io_matchBytes_1332(matchBytes[1332]),
.io_matchBytes_1333(matchBytes[1333]),
.io_matchBytes_1334(matchBytes[1334]),
.io_matchBytes_1335(matchBytes[1335]),
.io_matchBytes_1336(matchBytes[1336]),
.io_matchBytes_1337(matchBytes[1337]),
.io_matchBytes_1338(matchBytes[1338]),
.io_matchBytes_1339(matchBytes[1339]),
.io_matchBytes_1340(matchBytes[1340]),
.io_matchBytes_1341(matchBytes[1341]),
.io_matchBytes_1342(matchBytes[1342]),
.io_matchBytes_1343(matchBytes[1343]),
.io_matchBytes_1344(matchBytes[1344]),
.io_matchBytes_1345(matchBytes[1345]),
.io_matchBytes_1346(matchBytes[1346]),
.io_matchBytes_1347(matchBytes[1347]),
.io_matchBytes_1348(matchBytes[1348]),
.io_matchBytes_1349(matchBytes[1349]),
.io_matchBytes_1350(matchBytes[1350]),
.io_matchBytes_1351(matchBytes[1351]),
.io_matchBytes_1352(matchBytes[1352]),
.io_matchBytes_1353(matchBytes[1353]),
.io_matchBytes_1354(matchBytes[1354]),
.io_matchBytes_1355(matchBytes[1355]),
.io_matchBytes_1356(matchBytes[1356]),
.io_matchBytes_1357(matchBytes[1357]),
.io_matchBytes_1358(matchBytes[1358]),
.io_matchBytes_1359(matchBytes[1359]),
.io_matchBytes_1360(matchBytes[1360]),
.io_matchBytes_1361(matchBytes[1361]),
.io_matchBytes_1362(matchBytes[1362]),
.io_matchBytes_1363(matchBytes[1363]),
.io_matchBytes_1364(matchBytes[1364]),
.io_matchBytes_1365(matchBytes[1365]),
.io_matchBytes_1366(matchBytes[1366]),
.io_matchBytes_1367(matchBytes[1367]),
.io_matchBytes_1368(matchBytes[1368]),
.io_matchBytes_1369(matchBytes[1369]),
.io_matchBytes_1370(matchBytes[1370]),
.io_matchBytes_1371(matchBytes[1371]),
.io_matchBytes_1372(matchBytes[1372]),
.io_matchBytes_1373(matchBytes[1373]),
.io_matchBytes_1374(matchBytes[1374]),
.io_matchBytes_1375(matchBytes[1375]),
.io_matchBytes_1376(matchBytes[1376]),
.io_matchBytes_1377(matchBytes[1377]),
.io_matchBytes_1378(matchBytes[1378]),
.io_matchBytes_1379(matchBytes[1379]),
.io_matchBytes_1380(matchBytes[1380]),
.io_matchBytes_1381(matchBytes[1381]),
.io_matchBytes_1382(matchBytes[1382]),
.io_matchBytes_1383(matchBytes[1383]),
.io_matchBytes_1384(matchBytes[1384]),
.io_matchBytes_1385(matchBytes[1385]),
.io_matchBytes_1386(matchBytes[1386]),
.io_matchBytes_1387(matchBytes[1387]),
.io_matchBytes_1388(matchBytes[1388]),
.io_matchBytes_1389(matchBytes[1389]),
.io_matchBytes_1390(matchBytes[1390]),
.io_matchBytes_1391(matchBytes[1391]),
.io_matchBytes_1392(matchBytes[1392]),
.io_matchBytes_1393(matchBytes[1393]),
.io_matchBytes_1394(matchBytes[1394]),
.io_matchBytes_1395(matchBytes[1395]),
.io_matchBytes_1396(matchBytes[1396]),
.io_matchBytes_1397(matchBytes[1397]),
.io_matchBytes_1398(matchBytes[1398]),
.io_matchBytes_1399(matchBytes[1399]),
.io_matchBytes_1400(matchBytes[1400]),
.io_matchBytes_1401(matchBytes[1401]),
.io_matchBytes_1402(matchBytes[1402]),
.io_matchBytes_1403(matchBytes[1403]),
.io_matchBytes_1404(matchBytes[1404]),
.io_matchBytes_1405(matchBytes[1405]),
.io_matchBytes_1406(matchBytes[1406]),
.io_matchBytes_1407(matchBytes[1407]),
.io_matchBytes_1408(matchBytes[1408]),
.io_matchBytes_1409(matchBytes[1409]),
.io_matchBytes_1410(matchBytes[1410]),
.io_matchBytes_1411(matchBytes[1411]),
.io_matchBytes_1412(matchBytes[1412]),
.io_matchBytes_1413(matchBytes[1413]),
.io_matchBytes_1414(matchBytes[1414]),
.io_matchBytes_1415(matchBytes[1415]),
.io_matchBytes_1416(matchBytes[1416]),
.io_matchBytes_1417(matchBytes[1417]),
.io_matchBytes_1418(matchBytes[1418]),
.io_matchBytes_1419(matchBytes[1419]),
.io_matchBytes_1420(matchBytes[1420]),
.io_matchBytes_1421(matchBytes[1421]),
.io_matchBytes_1422(matchBytes[1422]),
.io_matchBytes_1423(matchBytes[1423]),
.io_matchBytes_1424(matchBytes[1424]),
.io_matchBytes_1425(matchBytes[1425]),
.io_matchBytes_1426(matchBytes[1426]),
.io_matchBytes_1427(matchBytes[1427]),
.io_matchBytes_1428(matchBytes[1428]),
.io_matchBytes_1429(matchBytes[1429]),
.io_matchBytes_1430(matchBytes[1430]),
.io_matchBytes_1431(matchBytes[1431]),
.io_matchBytes_1432(matchBytes[1432]),
.io_matchBytes_1433(matchBytes[1433]),
.io_matchBytes_1434(matchBytes[1434]),
.io_matchBytes_1435(matchBytes[1435]),
.io_matchBytes_1436(matchBytes[1436]),
.io_matchBytes_1437(matchBytes[1437]),
.io_matchBytes_1438(matchBytes[1438]),
.io_matchBytes_1439(matchBytes[1439]),
.io_matchBytes_1440(matchBytes[1440]),
.io_matchBytes_1441(matchBytes[1441]),
.io_matchBytes_1442(matchBytes[1442]),
.io_matchBytes_1443(matchBytes[1443]),
.io_matchBytes_1444(matchBytes[1444]),
.io_matchBytes_1445(matchBytes[1445]),
.io_matchBytes_1446(matchBytes[1446]),
.io_matchBytes_1447(matchBytes[1447]),
.io_matchBytes_1448(matchBytes[1448]),
.io_matchBytes_1449(matchBytes[1449]),
.io_matchBytes_1450(matchBytes[1450]),
.io_matchBytes_1451(matchBytes[1451]),
.io_matchBytes_1452(matchBytes[1452]),
.io_matchBytes_1453(matchBytes[1453]),
.io_matchBytes_1454(matchBytes[1454]),
.io_matchBytes_1455(matchBytes[1455]),
.io_matchBytes_1456(matchBytes[1456]),
.io_matchBytes_1457(matchBytes[1457]),
.io_matchBytes_1458(matchBytes[1458]),
.io_matchBytes_1459(matchBytes[1459]),
.io_matchBytes_1460(matchBytes[1460]),
.io_matchBytes_1461(matchBytes[1461]),
.io_matchBytes_1462(matchBytes[1462]),
.io_matchBytes_1463(matchBytes[1463]),
.io_matchBytes_1464(matchBytes[1464]),
.io_matchBytes_1465(matchBytes[1465]),
.io_matchBytes_1466(matchBytes[1466]),
.io_matchBytes_1467(matchBytes[1467]),
.io_matchBytes_1468(matchBytes[1468]),
.io_matchBytes_1469(matchBytes[1469]),
.io_matchBytes_1470(matchBytes[1470]),
.io_matchBytes_1471(matchBytes[1471]),
.io_matchBytes_1472(matchBytes[1472]),
.io_matchBytes_1473(matchBytes[1473]),
.io_matchBytes_1474(matchBytes[1474]),
.io_matchBytes_1475(matchBytes[1475]),
.io_matchBytes_1476(matchBytes[1476]),
.io_matchBytes_1477(matchBytes[1477]),
.io_matchBytes_1478(matchBytes[1478]),
.io_matchBytes_1479(matchBytes[1479]),
.io_matchBytes_1480(matchBytes[1480]),
.io_matchBytes_1481(matchBytes[1481]),
.io_matchBytes_1482(matchBytes[1482]),
.io_matchBytes_1483(matchBytes[1483]),
.io_matchBytes_1484(matchBytes[1484]),
.io_matchBytes_1485(matchBytes[1485]),
.io_matchBytes_1486(matchBytes[1486]),
.io_matchBytes_1487(matchBytes[1487]),
.io_matchBytes_1488(matchBytes[1488]),
.io_matchBytes_1489(matchBytes[1489]),
.io_matchBytes_1490(matchBytes[1490]),
.io_matchBytes_1491(matchBytes[1491]),
.io_matchBytes_1492(matchBytes[1492]),
.io_matchBytes_1493(matchBytes[1493]),
.io_matchBytes_1494(matchBytes[1494]),
.io_matchBytes_1495(matchBytes[1495]),
.io_matchBytes_1496(matchBytes[1496]),
.io_matchBytes_1497(matchBytes[1497]),
.io_matchBytes_1498(matchBytes[1498]),
.io_matchBytes_1499(matchBytes[1499]),
.io_matchBytes_1500(matchBytes[1500]),
.io_matchBytes_1501(matchBytes[1501]),
.io_matchBytes_1502(matchBytes[1502]),
.io_matchBytes_1503(matchBytes[1503]),
.io_matchBytes_1504(matchBytes[1504]),
.io_matchBytes_1505(matchBytes[1505]),
.io_matchBytes_1506(matchBytes[1506]),
.io_matchBytes_1507(matchBytes[1507]),
.io_matchBytes_1508(matchBytes[1508]),
.io_matchBytes_1509(matchBytes[1509]),
.io_matchBytes_1510(matchBytes[1510]),
.io_matchBytes_1511(matchBytes[1511]),
.io_matchBytes_1512(matchBytes[1512]),
.io_matchBytes_1513(matchBytes[1513]),
.io_matchBytes_1514(matchBytes[1514]),
.io_matchBytes_1515(matchBytes[1515]),
.io_matchBytes_1516(matchBytes[1516]),
.io_matchBytes_1517(matchBytes[1517]),
.io_matchBytes_1518(matchBytes[1518]),
.io_matchBytes_1519(matchBytes[1519]),
.io_matchBytes_1520(matchBytes[1520]),
.io_matchBytes_1521(matchBytes[1521]),
.io_matchBytes_1522(matchBytes[1522]),
.io_matchBytes_1523(matchBytes[1523]),
.io_matchBytes_1524(matchBytes[1524]),
.io_matchBytes_1525(matchBytes[1525]),
.io_matchBytes_1526(matchBytes[1526]),
.io_matchBytes_1527(matchBytes[1527]),
.io_matchBytes_1528(matchBytes[1528]),
.io_matchBytes_1529(matchBytes[1529]),
.io_matchBytes_1530(matchBytes[1530]),
.io_matchBytes_1531(matchBytes[1531]),
.io_matchBytes_1532(matchBytes[1532]),
.io_matchBytes_1533(matchBytes[1533]),
.io_matchBytes_1534(matchBytes[1534]),
.io_matchBytes_1535(matchBytes[1535]),
.io_matchBytes_1536(matchBytes[1536]),
.io_matchBytes_1537(matchBytes[1537]),
.io_matchBytes_1538(matchBytes[1538]),
.io_matchBytes_1539(matchBytes[1539]),
.io_matchBytes_1540(matchBytes[1540]),
.io_matchBytes_1541(matchBytes[1541]),
.io_matchBytes_1542(matchBytes[1542]),
.io_matchBytes_1543(matchBytes[1543]),
.io_matchBytes_1544(matchBytes[1544]),
.io_matchBytes_1545(matchBytes[1545]),
.io_matchBytes_1546(matchBytes[1546]),
.io_matchBytes_1547(matchBytes[1547]),
.io_matchBytes_1548(matchBytes[1548]),
.io_matchBytes_1549(matchBytes[1549]),
.io_matchBytes_1550(matchBytes[1550]),
.io_matchBytes_1551(matchBytes[1551]),
.io_matchBytes_1552(matchBytes[1552]),
.io_matchBytes_1553(matchBytes[1553]),
.io_matchBytes_1554(matchBytes[1554]),
.io_matchBytes_1555(matchBytes[1555]),
.io_matchBytes_1556(matchBytes[1556]),
.io_matchBytes_1557(matchBytes[1557]),
.io_matchBytes_1558(matchBytes[1558]),
.io_matchBytes_1559(matchBytes[1559]),
.io_matchBytes_1560(matchBytes[1560]),
.io_matchBytes_1561(matchBytes[1561]),
.io_matchBytes_1562(matchBytes[1562]),
.io_matchBytes_1563(matchBytes[1563]),
.io_matchBytes_1564(matchBytes[1564]),
.io_matchBytes_1565(matchBytes[1565]),
.io_matchBytes_1566(matchBytes[1566]),
.io_matchBytes_1567(matchBytes[1567]),
.io_matchBytes_1568(matchBytes[1568]),
.io_matchBytes_1569(matchBytes[1569]),
.io_matchBytes_1570(matchBytes[1570]),
.io_matchBytes_1571(matchBytes[1571]),
.io_matchBytes_1572(matchBytes[1572]),
.io_matchBytes_1573(matchBytes[1573]),
.io_matchBytes_1574(matchBytes[1574]),
.io_matchBytes_1575(matchBytes[1575]),
.io_matchBytes_1576(matchBytes[1576]),
.io_matchBytes_1577(matchBytes[1577]),
.io_matchBytes_1578(matchBytes[1578]),
.io_matchBytes_1579(matchBytes[1579]),
.io_matchBytes_1580(matchBytes[1580]),
.io_matchBytes_1581(matchBytes[1581]),
.io_matchBytes_1582(matchBytes[1582]),
.io_matchBytes_1583(matchBytes[1583]),
.io_matchBytes_1584(matchBytes[1584]),
.io_matchBytes_1585(matchBytes[1585]),
.io_matchBytes_1586(matchBytes[1586]),
.io_matchBytes_1587(matchBytes[1587]),
.io_matchBytes_1588(matchBytes[1588]),
.io_matchBytes_1589(matchBytes[1589]),
.io_matchBytes_1590(matchBytes[1590]),
.io_matchBytes_1591(matchBytes[1591]),
.io_matchBytes_1592(matchBytes[1592]),
.io_matchBytes_1593(matchBytes[1593]),
.io_matchBytes_1594(matchBytes[1594]),
.io_matchBytes_1595(matchBytes[1595]),
.io_matchBytes_1596(matchBytes[1596]),
.io_matchBytes_1597(matchBytes[1597]),
.io_matchBytes_1598(matchBytes[1598]),
.io_matchBytes_1599(matchBytes[1599]),
.io_matchBytes_1600(matchBytes[1600]),
.io_matchBytes_1601(matchBytes[1601]),
.io_matchBytes_1602(matchBytes[1602]),
.io_matchBytes_1603(matchBytes[1603]),
.io_matchBytes_1604(matchBytes[1604]),
.io_matchBytes_1605(matchBytes[1605]),
.io_matchBytes_1606(matchBytes[1606]),
.io_matchBytes_1607(matchBytes[1607]),
.io_matchBytes_1608(matchBytes[1608]),
.io_matchBytes_1609(matchBytes[1609]),
.io_matchBytes_1610(matchBytes[1610]),
.io_matchBytes_1611(matchBytes[1611]),
.io_matchBytes_1612(matchBytes[1612]),
.io_matchBytes_1613(matchBytes[1613]),
.io_matchBytes_1614(matchBytes[1614]),
.io_matchBytes_1615(matchBytes[1615]),
.io_matchBytes_1616(matchBytes[1616]),
.io_matchBytes_1617(matchBytes[1617]),
.io_matchBytes_1618(matchBytes[1618]),
.io_matchBytes_1619(matchBytes[1619]),
.io_matchBytes_1620(matchBytes[1620]),
.io_matchBytes_1621(matchBytes[1621]),
.io_matchBytes_1622(matchBytes[1622]),
.io_matchBytes_1623(matchBytes[1623]),
.io_matchBytes_1624(matchBytes[1624]),
.io_matchBytes_1625(matchBytes[1625]),
.io_matchBytes_1626(matchBytes[1626]),
.io_matchBytes_1627(matchBytes[1627]),
.io_matchBytes_1628(matchBytes[1628]),
.io_matchBytes_1629(matchBytes[1629]),
.io_matchBytes_1630(matchBytes[1630]),
.io_matchBytes_1631(matchBytes[1631]),
.io_matchBytes_1632(matchBytes[1632]),
.io_matchBytes_1633(matchBytes[1633]),
.io_matchBytes_1634(matchBytes[1634]),
.io_matchBytes_1635(matchBytes[1635]),
.io_matchBytes_1636(matchBytes[1636]),
.io_matchBytes_1637(matchBytes[1637]),
.io_matchBytes_1638(matchBytes[1638]),
.io_matchBytes_1639(matchBytes[1639]),
.io_matchBytes_1640(matchBytes[1640]),
.io_matchBytes_1641(matchBytes[1641]),
.io_matchBytes_1642(matchBytes[1642]),
.io_matchBytes_1643(matchBytes[1643]),
.io_matchBytes_1644(matchBytes[1644]),
.io_matchBytes_1645(matchBytes[1645]),
.io_matchBytes_1646(matchBytes[1646]),
.io_matchBytes_1647(matchBytes[1647]),
.io_matchBytes_1648(matchBytes[1648]),
.io_matchBytes_1649(matchBytes[1649]),
.io_matchBytes_1650(matchBytes[1650]),
.io_matchBytes_1651(matchBytes[1651]),
.io_matchBytes_1652(matchBytes[1652]),
.io_matchBytes_1653(matchBytes[1653]),
.io_matchBytes_1654(matchBytes[1654]),
.io_matchBytes_1655(matchBytes[1655]),
.io_matchBytes_1656(matchBytes[1656]),
.io_matchBytes_1657(matchBytes[1657]),
.io_matchBytes_1658(matchBytes[1658]),
.io_matchBytes_1659(matchBytes[1659]),
.io_matchBytes_1660(matchBytes[1660]),
.io_matchBytes_1661(matchBytes[1661]),
.io_matchBytes_1662(matchBytes[1662]),
.io_matchBytes_1663(matchBytes[1663]),
.io_matchBytes_1664(matchBytes[1664]),
.io_matchBytes_1665(matchBytes[1665]),
.io_matchBytes_1666(matchBytes[1666]),
.io_matchBytes_1667(matchBytes[1667]),
.io_matchBytes_1668(matchBytes[1668]),
.io_matchBytes_1669(matchBytes[1669]),
.io_matchBytes_1670(matchBytes[1670]),
.io_matchBytes_1671(matchBytes[1671]),
.io_matchBytes_1672(matchBytes[1672]),
.io_matchBytes_1673(matchBytes[1673]),
.io_matchBytes_1674(matchBytes[1674]),
.io_matchBytes_1675(matchBytes[1675]),
.io_matchBytes_1676(matchBytes[1676]),
.io_matchBytes_1677(matchBytes[1677]),
.io_matchBytes_1678(matchBytes[1678]),
.io_matchBytes_1679(matchBytes[1679]),
.io_matchBytes_1680(matchBytes[1680]),
.io_matchBytes_1681(matchBytes[1681]),
.io_matchBytes_1682(matchBytes[1682]),
.io_matchBytes_1683(matchBytes[1683]),
.io_matchBytes_1684(matchBytes[1684]),
.io_matchBytes_1685(matchBytes[1685]),
.io_matchBytes_1686(matchBytes[1686]),
.io_matchBytes_1687(matchBytes[1687]),
.io_matchBytes_1688(matchBytes[1688]),
.io_matchBytes_1689(matchBytes[1689]),
.io_matchBytes_1690(matchBytes[1690]),
.io_matchBytes_1691(matchBytes[1691]),
.io_matchBytes_1692(matchBytes[1692]),
.io_matchBytes_1693(matchBytes[1693]),
.io_matchBytes_1694(matchBytes[1694]),
.io_matchBytes_1695(matchBytes[1695]),
.io_matchBytes_1696(matchBytes[1696]),
.io_matchBytes_1697(matchBytes[1697]),
.io_matchBytes_1698(matchBytes[1698]),
.io_matchBytes_1699(matchBytes[1699]),
.io_matchBytes_1700(matchBytes[1700]),
.io_matchBytes_1701(matchBytes[1701]),
.io_matchBytes_1702(matchBytes[1702]),
.io_matchBytes_1703(matchBytes[1703]),
.io_matchBytes_1704(matchBytes[1704]),
.io_matchBytes_1705(matchBytes[1705]),
.io_matchBytes_1706(matchBytes[1706]),
.io_matchBytes_1707(matchBytes[1707]),
.io_matchBytes_1708(matchBytes[1708]),
.io_matchBytes_1709(matchBytes[1709]),
.io_matchBytes_1710(matchBytes[1710]),
.io_matchBytes_1711(matchBytes[1711]),
.io_matchBytes_1712(matchBytes[1712]),
.io_matchBytes_1713(matchBytes[1713]),
.io_matchBytes_1714(matchBytes[1714]),
.io_matchBytes_1715(matchBytes[1715]),
.io_matchBytes_1716(matchBytes[1716]),
.io_matchBytes_1717(matchBytes[1717]),
.io_matchBytes_1718(matchBytes[1718]),
.io_matchBytes_1719(matchBytes[1719]),
.io_matchBytes_1720(matchBytes[1720]),
.io_matchBytes_1721(matchBytes[1721]),
.io_matchBytes_1722(matchBytes[1722]),
.io_matchBytes_1723(matchBytes[1723]),
.io_matchBytes_1724(matchBytes[1724]),
.io_matchBytes_1725(matchBytes[1725]),
.io_matchBytes_1726(matchBytes[1726]),
.io_matchBytes_1727(matchBytes[1727]),
.io_matchBytes_1728(matchBytes[1728]),
.io_matchBytes_1729(matchBytes[1729]),
.io_matchBytes_1730(matchBytes[1730]),
.io_matchBytes_1731(matchBytes[1731]),
.io_matchBytes_1732(matchBytes[1732]),
.io_matchBytes_1733(matchBytes[1733]),
.io_matchBytes_1734(matchBytes[1734]),
.io_matchBytes_1735(matchBytes[1735]),
.io_matchBytes_1736(matchBytes[1736]),
.io_matchBytes_1737(matchBytes[1737]),
.io_matchBytes_1738(matchBytes[1738]),
.io_matchBytes_1739(matchBytes[1739]),
.io_matchBytes_1740(matchBytes[1740]),
.io_matchBytes_1741(matchBytes[1741]),
.io_matchBytes_1742(matchBytes[1742]),
.io_matchBytes_1743(matchBytes[1743]),
.io_matchBytes_1744(matchBytes[1744]),
.io_matchBytes_1745(matchBytes[1745]),
.io_matchBytes_1746(matchBytes[1746]),
.io_matchBytes_1747(matchBytes[1747]),
.io_matchBytes_1748(matchBytes[1748]),
.io_matchBytes_1749(matchBytes[1749]),
.io_matchBytes_1750(matchBytes[1750]),
.io_matchBytes_1751(matchBytes[1751]),
.io_matchBytes_1752(matchBytes[1752]),
.io_matchBytes_1753(matchBytes[1753]),
.io_matchBytes_1754(matchBytes[1754]),
.io_matchBytes_1755(matchBytes[1755]),
.io_matchBytes_1756(matchBytes[1756]),
.io_matchBytes_1757(matchBytes[1757]),
.io_matchBytes_1758(matchBytes[1758]),
.io_matchBytes_1759(matchBytes[1759]),
.io_matchBytes_1760(matchBytes[1760]),
.io_matchBytes_1761(matchBytes[1761]),
.io_matchBytes_1762(matchBytes[1762]),
.io_matchBytes_1763(matchBytes[1763]),
.io_matchBytes_1764(matchBytes[1764]),
.io_matchBytes_1765(matchBytes[1765]),
.io_matchBytes_1766(matchBytes[1766]),
.io_matchBytes_1767(matchBytes[1767]),
.io_matchBytes_1768(matchBytes[1768]),
.io_matchBytes_1769(matchBytes[1769]),
.io_matchBytes_1770(matchBytes[1770]),
.io_matchBytes_1771(matchBytes[1771]),
.io_matchBytes_1772(matchBytes[1772]),
.io_matchBytes_1773(matchBytes[1773]),
.io_matchBytes_1774(matchBytes[1774]),
.io_matchBytes_1775(matchBytes[1775]),
.io_matchBytes_1776(matchBytes[1776]),
.io_matchBytes_1777(matchBytes[1777]),
.io_matchBytes_1778(matchBytes[1778]),
.io_matchBytes_1779(matchBytes[1779]),
.io_matchBytes_1780(matchBytes[1780]),
.io_matchBytes_1781(matchBytes[1781]),
.io_matchBytes_1782(matchBytes[1782]),
.io_matchBytes_1783(matchBytes[1783]),
.io_matchBytes_1784(matchBytes[1784]),
.io_matchBytes_1785(matchBytes[1785]),
.io_matchBytes_1786(matchBytes[1786]),
.io_matchBytes_1787(matchBytes[1787]),
.io_matchBytes_1788(matchBytes[1788]),
.io_matchBytes_1789(matchBytes[1789]),
.io_matchBytes_1790(matchBytes[1790]),
.io_matchBytes_1791(matchBytes[1791]),
.io_matchBytes_1792(matchBytes[1792]),
.io_matchBytes_1793(matchBytes[1793]),
.io_matchBytes_1794(matchBytes[1794]),
.io_matchBytes_1795(matchBytes[1795]),
.io_matchBytes_1796(matchBytes[1796]),
.io_matchBytes_1797(matchBytes[1797]),
.io_matchBytes_1798(matchBytes[1798]),
.io_matchBytes_1799(matchBytes[1799]),
.io_matchBytes_1800(matchBytes[1800]),
.io_matchBytes_1801(matchBytes[1801]),
.io_matchBytes_1802(matchBytes[1802]),
.io_matchBytes_1803(matchBytes[1803]),
.io_matchBytes_1804(matchBytes[1804]),
.io_matchBytes_1805(matchBytes[1805]),
.io_matchBytes_1806(matchBytes[1806]),
.io_matchBytes_1807(matchBytes[1807]),
.io_matchBytes_1808(matchBytes[1808]),
.io_matchBytes_1809(matchBytes[1809]),
.io_matchBytes_1810(matchBytes[1810]),
.io_matchBytes_1811(matchBytes[1811]),
.io_matchBytes_1812(matchBytes[1812]),
.io_matchBytes_1813(matchBytes[1813]),
.io_matchBytes_1814(matchBytes[1814]),
.io_matchBytes_1815(matchBytes[1815]),
.io_matchBytes_1816(matchBytes[1816]),
.io_matchBytes_1817(matchBytes[1817]),
.io_matchBytes_1818(matchBytes[1818]),
.io_matchBytes_1819(matchBytes[1819]),
.io_matchBytes_1820(matchBytes[1820]),
.io_matchBytes_1821(matchBytes[1821]),
.io_matchBytes_1822(matchBytes[1822]),
.io_matchBytes_1823(matchBytes[1823]),
.io_matchBytes_1824(matchBytes[1824]),
.io_matchBytes_1825(matchBytes[1825]),
.io_matchBytes_1826(matchBytes[1826]),
.io_matchBytes_1827(matchBytes[1827]),
.io_matchBytes_1828(matchBytes[1828]),
.io_matchBytes_1829(matchBytes[1829]),
.io_matchBytes_1830(matchBytes[1830]),
.io_matchBytes_1831(matchBytes[1831]),
.io_matchBytes_1832(matchBytes[1832]),
.io_matchBytes_1833(matchBytes[1833]),
.io_matchBytes_1834(matchBytes[1834]),
.io_matchBytes_1835(matchBytes[1835]),
.io_matchBytes_1836(matchBytes[1836]),
.io_matchBytes_1837(matchBytes[1837]),
.io_matchBytes_1838(matchBytes[1838]),
.io_matchBytes_1839(matchBytes[1839]),
.io_matchBytes_1840(matchBytes[1840]),
.io_matchBytes_1841(matchBytes[1841]),
.io_matchBytes_1842(matchBytes[1842]),
.io_matchBytes_1843(matchBytes[1843]),
.io_matchBytes_1844(matchBytes[1844]),
.io_matchBytes_1845(matchBytes[1845]),
.io_matchBytes_1846(matchBytes[1846]),
.io_matchBytes_1847(matchBytes[1847]),
.io_matchBytes_1848(matchBytes[1848]),
.io_matchBytes_1849(matchBytes[1849]),
.io_matchBytes_1850(matchBytes[1850]),
.io_matchBytes_1851(matchBytes[1851]),
.io_matchBytes_1852(matchBytes[1852]),
.io_matchBytes_1853(matchBytes[1853]),
.io_matchBytes_1854(matchBytes[1854]),
.io_matchBytes_1855(matchBytes[1855]),
.io_matchBytes_1856(matchBytes[1856]),
.io_matchBytes_1857(matchBytes[1857]),
.io_matchBytes_1858(matchBytes[1858]),
.io_matchBytes_1859(matchBytes[1859]),
.io_matchBytes_1860(matchBytes[1860]),
.io_matchBytes_1861(matchBytes[1861]),
.io_matchBytes_1862(matchBytes[1862]),
.io_matchBytes_1863(matchBytes[1863]),
.io_matchBytes_1864(matchBytes[1864]),
.io_matchBytes_1865(matchBytes[1865]),
.io_matchBytes_1866(matchBytes[1866]),
.io_matchBytes_1867(matchBytes[1867]),
.io_matchBytes_1868(matchBytes[1868]),
.io_matchBytes_1869(matchBytes[1869]),
.io_matchBytes_1870(matchBytes[1870]),
.io_matchBytes_1871(matchBytes[1871]),
.io_matchBytes_1872(matchBytes[1872]),
.io_matchBytes_1873(matchBytes[1873]),
.io_matchBytes_1874(matchBytes[1874]),
.io_matchBytes_1875(matchBytes[1875]),
.io_matchBytes_1876(matchBytes[1876]),
.io_matchBytes_1877(matchBytes[1877]),
.io_matchBytes_1878(matchBytes[1878]),
.io_matchBytes_1879(matchBytes[1879]),
.io_matchBytes_1880(matchBytes[1880]),
.io_matchBytes_1881(matchBytes[1881]),
.io_matchBytes_1882(matchBytes[1882]),
.io_matchBytes_1883(matchBytes[1883]),
.io_matchBytes_1884(matchBytes[1884]),
.io_matchBytes_1885(matchBytes[1885]),
.io_matchBytes_1886(matchBytes[1886]),
.io_matchBytes_1887(matchBytes[1887]),
.io_matchBytes_1888(matchBytes[1888]),
.io_matchBytes_1889(matchBytes[1889]),
.io_matchBytes_1890(matchBytes[1890]),
.io_matchBytes_1891(matchBytes[1891]),
.io_matchBytes_1892(matchBytes[1892]),
.io_matchBytes_1893(matchBytes[1893]),
.io_matchBytes_1894(matchBytes[1894]),
.io_matchBytes_1895(matchBytes[1895]),
.io_matchBytes_1896(matchBytes[1896]),
.io_matchBytes_1897(matchBytes[1897]),
.io_matchBytes_1898(matchBytes[1898]),
.io_matchBytes_1899(matchBytes[1899]),
.io_matchBytes_1900(matchBytes[1900]),
.io_matchBytes_1901(matchBytes[1901]),
.io_matchBytes_1902(matchBytes[1902]),
.io_matchBytes_1903(matchBytes[1903]),
.io_matchBytes_1904(matchBytes[1904]),
.io_matchBytes_1905(matchBytes[1905]),
.io_matchBytes_1906(matchBytes[1906]),
.io_matchBytes_1907(matchBytes[1907]),
.io_matchBytes_1908(matchBytes[1908]),
.io_matchBytes_1909(matchBytes[1909]),
.io_matchBytes_1910(matchBytes[1910]),
.io_matchBytes_1911(matchBytes[1911]),
.io_matchBytes_1912(matchBytes[1912]),
.io_matchBytes_1913(matchBytes[1913]),
.io_matchBytes_1914(matchBytes[1914]),
.io_matchBytes_1915(matchBytes[1915]),
.io_matchBytes_1916(matchBytes[1916]),
.io_matchBytes_1917(matchBytes[1917]),
.io_matchBytes_1918(matchBytes[1918]),
.io_matchBytes_1919(matchBytes[1919]),
.io_matchBytes_1920(matchBytes[1920]),
.io_matchBytes_1921(matchBytes[1921]),
.io_matchBytes_1922(matchBytes[1922]),
.io_matchBytes_1923(matchBytes[1923]),
.io_matchBytes_1924(matchBytes[1924]),
.io_matchBytes_1925(matchBytes[1925]),
.io_matchBytes_1926(matchBytes[1926]),
.io_matchBytes_1927(matchBytes[1927]),
.io_matchBytes_1928(matchBytes[1928]),
.io_matchBytes_1929(matchBytes[1929]),
.io_matchBytes_1930(matchBytes[1930]),
.io_matchBytes_1931(matchBytes[1931]),
.io_matchBytes_1932(matchBytes[1932]),
.io_matchBytes_1933(matchBytes[1933]),
.io_matchBytes_1934(matchBytes[1934]),
.io_matchBytes_1935(matchBytes[1935]),
.io_matchBytes_1936(matchBytes[1936]),
.io_matchBytes_1937(matchBytes[1937]),
.io_matchBytes_1938(matchBytes[1938]),
.io_matchBytes_1939(matchBytes[1939]),
.io_matchBytes_1940(matchBytes[1940]),
.io_matchBytes_1941(matchBytes[1941]),
.io_matchBytes_1942(matchBytes[1942]),
.io_matchBytes_1943(matchBytes[1943]),
.io_matchBytes_1944(matchBytes[1944]),
.io_matchBytes_1945(matchBytes[1945]),
.io_matchBytes_1946(matchBytes[1946]),
.io_matchBytes_1947(matchBytes[1947]),
.io_matchBytes_1948(matchBytes[1948]),
.io_matchBytes_1949(matchBytes[1949]),
.io_matchBytes_1950(matchBytes[1950]),
.io_matchBytes_1951(matchBytes[1951]),
.io_matchBytes_1952(matchBytes[1952]),
.io_matchBytes_1953(matchBytes[1953]),
.io_matchBytes_1954(matchBytes[1954]),
.io_matchBytes_1955(matchBytes[1955]),
.io_matchBytes_1956(matchBytes[1956]),
.io_matchBytes_1957(matchBytes[1957]),
.io_matchBytes_1958(matchBytes[1958]),
.io_matchBytes_1959(matchBytes[1959]),
.io_matchBytes_1960(matchBytes[1960]),
.io_matchBytes_1961(matchBytes[1961]),
.io_matchBytes_1962(matchBytes[1962]),
.io_matchBytes_1963(matchBytes[1963]),
.io_matchBytes_1964(matchBytes[1964]),
.io_matchBytes_1965(matchBytes[1965]),
.io_matchBytes_1966(matchBytes[1966]),
.io_matchBytes_1967(matchBytes[1967]),
.io_matchBytes_1968(matchBytes[1968]),
.io_matchBytes_1969(matchBytes[1969]),
.io_matchBytes_1970(matchBytes[1970]),
.io_matchBytes_1971(matchBytes[1971]),
.io_matchBytes_1972(matchBytes[1972]),
.io_matchBytes_1973(matchBytes[1973]),
.io_matchBytes_1974(matchBytes[1974]),
.io_matchBytes_1975(matchBytes[1975]),
.io_matchBytes_1976(matchBytes[1976]),
.io_matchBytes_1977(matchBytes[1977]),
.io_matchBytes_1978(matchBytes[1978]),
.io_matchBytes_1979(matchBytes[1979]),
.io_matchBytes_1980(matchBytes[1980]),
.io_matchBytes_1981(matchBytes[1981]),
.io_matchBytes_1982(matchBytes[1982]),
.io_matchBytes_1983(matchBytes[1983]),
.io_matchBytes_1984(matchBytes[1984]),
.io_matchBytes_1985(matchBytes[1985]),
.io_matchBytes_1986(matchBytes[1986]),
.io_matchBytes_1987(matchBytes[1987]),
.io_matchBytes_1988(matchBytes[1988]),
.io_matchBytes_1989(matchBytes[1989]),
.io_matchBytes_1990(matchBytes[1990]),
.io_matchBytes_1991(matchBytes[1991]),
.io_matchBytes_1992(matchBytes[1992]),
.io_matchBytes_1993(matchBytes[1993]),
.io_matchBytes_1994(matchBytes[1994]),
.io_matchBytes_1995(matchBytes[1995]),
.io_matchBytes_1996(matchBytes[1996]),
.io_matchBytes_1997(matchBytes[1997]),
.io_matchBytes_1998(matchBytes[1998]),
.io_matchBytes_1999(matchBytes[1999]),
.io_matchBytes_2000(matchBytes[2000]),
.io_matchBytes_2001(matchBytes[2001]),
.io_matchBytes_2002(matchBytes[2002]),
.io_matchBytes_2003(matchBytes[2003]),
.io_matchBytes_2004(matchBytes[2004]),
.io_matchBytes_2005(matchBytes[2005]),
.io_matchBytes_2006(matchBytes[2006]),
.io_matchBytes_2007(matchBytes[2007]),
.io_matchBytes_2008(matchBytes[2008]),
.io_matchBytes_2009(matchBytes[2009]),
.io_matchBytes_2010(matchBytes[2010]),
.io_matchBytes_2011(matchBytes[2011]),
.io_matchBytes_2012(matchBytes[2012]),
.io_matchBytes_2013(matchBytes[2013]),
.io_matchBytes_2014(matchBytes[2014]),
.io_matchBytes_2015(matchBytes[2015]),
.io_matchBytes_2016(matchBytes[2016]),
.io_matchBytes_2017(matchBytes[2017]),
.io_matchBytes_2018(matchBytes[2018]),
.io_matchBytes_2019(matchBytes[2019]),
.io_matchBytes_2020(matchBytes[2020]),
.io_matchBytes_2021(matchBytes[2021]),
.io_matchBytes_2022(matchBytes[2022]),
.io_matchBytes_2023(matchBytes[2023]),
.io_matchBytes_2024(matchBytes[2024]),
.io_matchBytes_2025(matchBytes[2025]),
.io_matchBytes_2026(matchBytes[2026]),
.io_matchBytes_2027(matchBytes[2027]),
.io_matchBytes_2028(matchBytes[2028]),
.io_matchBytes_2029(matchBytes[2029]),
.io_matchBytes_2030(matchBytes[2030]),
.io_matchBytes_2031(matchBytes[2031]),
.io_matchBytes_2032(matchBytes[2032]),
.io_matchBytes_2033(matchBytes[2033]),
.io_matchBytes_2034(matchBytes[2034]),
.io_matchBytes_2035(matchBytes[2035]),
.io_matchBytes_2036(matchBytes[2036]),
.io_matchBytes_2037(matchBytes[2037]),
.io_matchBytes_2038(matchBytes[2038]),
.io_matchBytes_2039(matchBytes[2039]),
.io_matchBytes_2040(matchBytes[2040]),
.io_matchBytes_2041(matchBytes[2041]),
.io_matchBytes_2042(matchBytes[2042]),
.io_matchBytes_2043(matchBytes[2043]),
.io_matchBytes_2044(matchBytes[2044]),
.io_matchBytes_2045(matchBytes[2045]),
.io_matchBytes_2046(matchBytes[2046]),
.io_matchBytes_2047(matchBytes[2047]),
.io_matchBytes_2048(matchBytes[2048]),
.io_matchBytes_2049(matchBytes[2049]),
.io_matchBytes_2050(matchBytes[2050]),
.io_matchBytes_2051(matchBytes[2051]),
.io_matchBytes_2052(matchBytes[2052]),
.io_matchBytes_2053(matchBytes[2053]),
.io_matchBytes_2054(matchBytes[2054]),
.io_matchBytes_2055(matchBytes[2055]),
.io_matchBytes_2056(matchBytes[2056]),
.io_matchBytes_2057(matchBytes[2057]),
.io_matchBytes_2058(matchBytes[2058]),
.io_matchBytes_2059(matchBytes[2059]),
.io_matchBytes_2060(matchBytes[2060]),
.io_matchBytes_2061(matchBytes[2061]),
.io_matchBytes_2062(matchBytes[2062]),
.io_matchBytes_2063(matchBytes[2063]),
.io_matchBytes_2064(matchBytes[2064]),
.io_matchBytes_2065(matchBytes[2065]),
.io_matchBytes_2066(matchBytes[2066]),
.io_matchBytes_2067(matchBytes[2067]),
.io_matchBytes_2068(matchBytes[2068]),
.io_matchBytes_2069(matchBytes[2069]),
.io_matchBytes_2070(matchBytes[2070]),
.io_matchBytes_2071(matchBytes[2071]),
.io_matchBytes_2072(matchBytes[2072]),
.io_matchBytes_2073(matchBytes[2073]),
.io_matchBytes_2074(matchBytes[2074]),
.io_matchBytes_2075(matchBytes[2075]),
.io_matchBytes_2076(matchBytes[2076]),
.io_matchBytes_2077(matchBytes[2077]),
.io_matchBytes_2078(matchBytes[2078]),
.io_matchBytes_2079(matchBytes[2079]),
.io_matchBytes_2080(matchBytes[2080]),
.io_matchBytes_2081(matchBytes[2081]),
.io_matchBytes_2082(matchBytes[2082]),
.io_matchBytes_2083(matchBytes[2083]),
.io_matchBytes_2084(matchBytes[2084]),
.io_matchBytes_2085(matchBytes[2085]),
.io_matchBytes_2086(matchBytes[2086]),
.io_matchBytes_2087(matchBytes[2087]),
.io_matchBytes_2088(matchBytes[2088]),
.io_matchBytes_2089(matchBytes[2089]),
.io_matchBytes_2090(matchBytes[2090]),
.io_matchBytes_2091(matchBytes[2091]),
.io_matchBytes_2092(matchBytes[2092]),
.io_matchBytes_2093(matchBytes[2093]),
.io_matchBytes_2094(matchBytes[2094]),
.io_matchBytes_2095(matchBytes[2095]),
.io_matchBytes_2096(matchBytes[2096]),
.io_matchBytes_2097(matchBytes[2097]),
.io_matchBytes_2098(matchBytes[2098]),
.io_matchBytes_2099(matchBytes[2099]),
.io_matchBytes_2100(matchBytes[2100]),
.io_matchBytes_2101(matchBytes[2101]),
.io_matchBytes_2102(matchBytes[2102]),
.io_matchBytes_2103(matchBytes[2103]),
.io_matchBytes_2104(matchBytes[2104]),
.io_matchBytes_2105(matchBytes[2105]),
.io_matchBytes_2106(matchBytes[2106]),
.io_matchBytes_2107(matchBytes[2107]),
.io_matchBytes_2108(matchBytes[2108]),
.io_matchBytes_2109(matchBytes[2109]),
.io_matchBytes_2110(matchBytes[2110]),
.io_matchBytes_2111(matchBytes[2111]),
.io_matchBytes_2112(matchBytes[2112]),
.io_matchBytes_2113(matchBytes[2113]),
.io_matchBytes_2114(matchBytes[2114]),
.io_matchBytes_2115(matchBytes[2115]),
.io_matchBytes_2116(matchBytes[2116]),
.io_matchBytes_2117(matchBytes[2117]),
.io_matchBytes_2118(matchBytes[2118]),
.io_matchBytes_2119(matchBytes[2119]),
.io_matchBytes_2120(matchBytes[2120]),
.io_matchBytes_2121(matchBytes[2121]),
.io_matchBytes_2122(matchBytes[2122]),
.io_matchBytes_2123(matchBytes[2123]),
.io_matchBytes_2124(matchBytes[2124]),
.io_matchBytes_2125(matchBytes[2125]),
.io_matchBytes_2126(matchBytes[2126]),
.io_matchBytes_2127(matchBytes[2127]),
.io_matchBytes_2128(matchBytes[2128]),
.io_matchBytes_2129(matchBytes[2129]),
.io_matchBytes_2130(matchBytes[2130]),
.io_matchBytes_2131(matchBytes[2131]),
.io_matchBytes_2132(matchBytes[2132]),
.io_matchBytes_2133(matchBytes[2133]),
.io_matchBytes_2134(matchBytes[2134]),
.io_matchBytes_2135(matchBytes[2135]),
.io_matchBytes_2136(matchBytes[2136]),
.io_matchBytes_2137(matchBytes[2137]),
.io_matchBytes_2138(matchBytes[2138]),
.io_matchBytes_2139(matchBytes[2139]),
.io_matchBytes_2140(matchBytes[2140]),
.io_matchBytes_2141(matchBytes[2141]),
.io_matchBytes_2142(matchBytes[2142]),
.io_matchBytes_2143(matchBytes[2143]),
.io_matchBytes_2144(matchBytes[2144]),
.io_matchBytes_2145(matchBytes[2145]),
.io_matchBytes_2146(matchBytes[2146]),
.io_matchBytes_2147(matchBytes[2147]),
.io_matchBytes_2148(matchBytes[2148]),
.io_matchBytes_2149(matchBytes[2149]),
.io_matchBytes_2150(matchBytes[2150]),
.io_matchBytes_2151(matchBytes[2151]),
.io_matchBytes_2152(matchBytes[2152]),
.io_matchBytes_2153(matchBytes[2153]),
.io_matchBytes_2154(matchBytes[2154]),
.io_matchBytes_2155(matchBytes[2155]),
.io_matchBytes_2156(matchBytes[2156]),
.io_matchBytes_2157(matchBytes[2157]),
.io_matchBytes_2158(matchBytes[2158]),
.io_matchBytes_2159(matchBytes[2159]),
.io_matchBytes_2160(matchBytes[2160]),
.io_matchBytes_2161(matchBytes[2161]),
.io_matchBytes_2162(matchBytes[2162]),
.io_matchBytes_2163(matchBytes[2163]),
.io_matchBytes_2164(matchBytes[2164]),
.io_matchBytes_2165(matchBytes[2165]),
.io_matchBytes_2166(matchBytes[2166]),
.io_matchBytes_2167(matchBytes[2167]),
.io_matchBytes_2168(matchBytes[2168]),
.io_matchBytes_2169(matchBytes[2169]),
.io_matchBytes_2170(matchBytes[2170]),
.io_matchBytes_2171(matchBytes[2171]),
.io_matchBytes_2172(matchBytes[2172]),
.io_matchBytes_2173(matchBytes[2173]),
.io_matchBytes_2174(matchBytes[2174]),
.io_matchBytes_2175(matchBytes[2175]),
.io_matchBytes_2176(matchBytes[2176]),
.io_matchBytes_2177(matchBytes[2177]),
.io_matchBytes_2178(matchBytes[2178]),
.io_matchBytes_2179(matchBytes[2179]),
.io_matchBytes_2180(matchBytes[2180]),
.io_matchBytes_2181(matchBytes[2181]),
.io_matchBytes_2182(matchBytes[2182]),
.io_matchBytes_2183(matchBytes[2183]),
.io_matchBytes_2184(matchBytes[2184]),
.io_matchBytes_2185(matchBytes[2185]),
.io_matchBytes_2186(matchBytes[2186]),
.io_matchBytes_2187(matchBytes[2187]),
.io_matchBytes_2188(matchBytes[2188]),
.io_matchBytes_2189(matchBytes[2189]),
.io_matchBytes_2190(matchBytes[2190]),
.io_matchBytes_2191(matchBytes[2191]),
.io_matchBytes_2192(matchBytes[2192]),
.io_matchBytes_2193(matchBytes[2193]),
.io_matchBytes_2194(matchBytes[2194]),
.io_matchBytes_2195(matchBytes[2195]),
.io_matchBytes_2196(matchBytes[2196]),
.io_matchBytes_2197(matchBytes[2197]),
.io_matchBytes_2198(matchBytes[2198]),
.io_matchBytes_2199(matchBytes[2199]),
.io_matchBytes_2200(matchBytes[2200]),
.io_matchBytes_2201(matchBytes[2201]),
.io_matchBytes_2202(matchBytes[2202]),
.io_matchBytes_2203(matchBytes[2203]),
.io_matchBytes_2204(matchBytes[2204]),
.io_matchBytes_2205(matchBytes[2205]),
.io_matchBytes_2206(matchBytes[2206]),
.io_matchBytes_2207(matchBytes[2207]),
.io_matchBytes_2208(matchBytes[2208]),
.io_matchBytes_2209(matchBytes[2209]),
.io_matchBytes_2210(matchBytes[2210]),
.io_matchBytes_2211(matchBytes[2211]),
.io_matchBytes_2212(matchBytes[2212]),
.io_matchBytes_2213(matchBytes[2213]),
.io_matchBytes_2214(matchBytes[2214]),
.io_matchBytes_2215(matchBytes[2215]),
.io_matchBytes_2216(matchBytes[2216]),
.io_matchBytes_2217(matchBytes[2217]),
.io_matchBytes_2218(matchBytes[2218]),
.io_matchBytes_2219(matchBytes[2219]),
.io_matchBytes_2220(matchBytes[2220]),
.io_matchBytes_2221(matchBytes[2221]),
.io_matchBytes_2222(matchBytes[2222]),
.io_matchBytes_2223(matchBytes[2223]),
.io_matchBytes_2224(matchBytes[2224]),
.io_matchBytes_2225(matchBytes[2225]),
.io_matchBytes_2226(matchBytes[2226]),
.io_matchBytes_2227(matchBytes[2227]),
.io_matchBytes_2228(matchBytes[2228]),
.io_matchBytes_2229(matchBytes[2229]),
.io_matchBytes_2230(matchBytes[2230]),
.io_matchBytes_2231(matchBytes[2231]),
.io_matchBytes_2232(matchBytes[2232]),
.io_matchBytes_2233(matchBytes[2233]),
.io_matchBytes_2234(matchBytes[2234]),
.io_matchBytes_2235(matchBytes[2235]),
.io_matchBytes_2236(matchBytes[2236]),
.io_matchBytes_2237(matchBytes[2237]),
.io_matchBytes_2238(matchBytes[2238]),
.io_matchBytes_2239(matchBytes[2239]),
.io_matchBytes_2240(matchBytes[2240]),
.io_matchBytes_2241(matchBytes[2241]),
.io_matchBytes_2242(matchBytes[2242]),
.io_matchBytes_2243(matchBytes[2243]),
.io_matchBytes_2244(matchBytes[2244]),
.io_matchBytes_2245(matchBytes[2245]),
.io_matchBytes_2246(matchBytes[2246]),
.io_matchBytes_2247(matchBytes[2247]),
.io_matchBytes_2248(matchBytes[2248]),
.io_matchBytes_2249(matchBytes[2249]),
.io_matchBytes_2250(matchBytes[2250]),
.io_matchBytes_2251(matchBytes[2251]),
.io_matchBytes_2252(matchBytes[2252]),
.io_matchBytes_2253(matchBytes[2253]),
.io_matchBytes_2254(matchBytes[2254]),
.io_matchBytes_2255(matchBytes[2255]),
.io_matchBytes_2256(matchBytes[2256]),
.io_matchBytes_2257(matchBytes[2257]),
.io_matchBytes_2258(matchBytes[2258]),
.io_matchBytes_2259(matchBytes[2259]),
.io_matchBytes_2260(matchBytes[2260]),
.io_matchBytes_2261(matchBytes[2261]),
.io_matchBytes_2262(matchBytes[2262]),
.io_matchBytes_2263(matchBytes[2263]),
.io_matchBytes_2264(matchBytes[2264]),
.io_matchBytes_2265(matchBytes[2265]),
.io_matchBytes_2266(matchBytes[2266]),
.io_matchBytes_2267(matchBytes[2267]),
.io_matchBytes_2268(matchBytes[2268]),
.io_matchBytes_2269(matchBytes[2269]),
.io_matchBytes_2270(matchBytes[2270]),
.io_matchBytes_2271(matchBytes[2271]),
.io_matchBytes_2272(matchBytes[2272]),
.io_matchBytes_2273(matchBytes[2273]),
.io_matchBytes_2274(matchBytes[2274]),
.io_matchBytes_2275(matchBytes[2275]),
.io_matchBytes_2276(matchBytes[2276]),
.io_matchBytes_2277(matchBytes[2277]),
.io_matchBytes_2278(matchBytes[2278]),
.io_matchBytes_2279(matchBytes[2279]),
.io_matchBytes_2280(matchBytes[2280]),
.io_matchBytes_2281(matchBytes[2281]),
.io_matchBytes_2282(matchBytes[2282]),
.io_matchBytes_2283(matchBytes[2283]),
.io_matchBytes_2284(matchBytes[2284]),
.io_matchBytes_2285(matchBytes[2285]),
.io_matchBytes_2286(matchBytes[2286]),
.io_matchBytes_2287(matchBytes[2287]),
.io_matchBytes_2288(matchBytes[2288]),
.io_matchBytes_2289(matchBytes[2289]),
.io_matchBytes_2290(matchBytes[2290]),
.io_matchBytes_2291(matchBytes[2291]),
.io_matchBytes_2292(matchBytes[2292]),
.io_matchBytes_2293(matchBytes[2293]),
.io_matchBytes_2294(matchBytes[2294]),
.io_matchBytes_2295(matchBytes[2295]),
.io_matchBytes_2296(matchBytes[2296]),
.io_matchBytes_2297(matchBytes[2297]),
.io_matchBytes_2298(matchBytes[2298]),
.io_matchBytes_2299(matchBytes[2299]),
.io_matchBytes_2300(matchBytes[2300]),
.io_matchBytes_2301(matchBytes[2301]),
.io_matchBytes_2302(matchBytes[2302]),
.io_matchBytes_2303(matchBytes[2303]),
.io_matchBytes_2304(matchBytes[2304]),
.io_matchBytes_2305(matchBytes[2305]),
.io_matchBytes_2306(matchBytes[2306]),
.io_matchBytes_2307(matchBytes[2307]),
.io_matchBytes_2308(matchBytes[2308]),
.io_matchBytes_2309(matchBytes[2309]),
.io_matchBytes_2310(matchBytes[2310]),
.io_matchBytes_2311(matchBytes[2311]),
.io_matchBytes_2312(matchBytes[2312]),
.io_matchBytes_2313(matchBytes[2313]),
.io_matchBytes_2314(matchBytes[2314]),
.io_matchBytes_2315(matchBytes[2315]),
.io_matchBytes_2316(matchBytes[2316]),
.io_matchBytes_2317(matchBytes[2317]),
.io_matchBytes_2318(matchBytes[2318]),
.io_matchBytes_2319(matchBytes[2319]),
.io_matchBytes_2320(matchBytes[2320]),
.io_matchBytes_2321(matchBytes[2321]),
.io_matchBytes_2322(matchBytes[2322]),
.io_matchBytes_2323(matchBytes[2323]),
.io_matchBytes_2324(matchBytes[2324]),
.io_matchBytes_2325(matchBytes[2325]),
.io_matchBytes_2326(matchBytes[2326]),
.io_matchBytes_2327(matchBytes[2327]),
.io_matchBytes_2328(matchBytes[2328]),
.io_matchBytes_2329(matchBytes[2329]),
.io_matchBytes_2330(matchBytes[2330]),
.io_matchBytes_2331(matchBytes[2331]),
.io_matchBytes_2332(matchBytes[2332]),
.io_matchBytes_2333(matchBytes[2333]),
.io_matchBytes_2334(matchBytes[2334]),
.io_matchBytes_2335(matchBytes[2335]),
.io_matchBytes_2336(matchBytes[2336]),
.io_matchBytes_2337(matchBytes[2337]),
.io_matchBytes_2338(matchBytes[2338]),
.io_matchBytes_2339(matchBytes[2339]),
.io_matchBytes_2340(matchBytes[2340]),
.io_matchBytes_2341(matchBytes[2341]),
.io_matchBytes_2342(matchBytes[2342]),
.io_matchBytes_2343(matchBytes[2343]),
.io_matchBytes_2344(matchBytes[2344]),
.io_matchBytes_2345(matchBytes[2345]),
.io_matchBytes_2346(matchBytes[2346]),
.io_matchBytes_2347(matchBytes[2347]),
.io_matchBytes_2348(matchBytes[2348]),
.io_matchBytes_2349(matchBytes[2349]),
.io_matchBytes_2350(matchBytes[2350]),
.io_matchBytes_2351(matchBytes[2351]),
.io_matchBytes_2352(matchBytes[2352]),
.io_matchBytes_2353(matchBytes[2353]),
.io_matchBytes_2354(matchBytes[2354]),
.io_matchBytes_2355(matchBytes[2355]),
.io_matchBytes_2356(matchBytes[2356]),
.io_matchBytes_2357(matchBytes[2357]),
.io_matchBytes_2358(matchBytes[2358]),
.io_matchBytes_2359(matchBytes[2359]),
.io_matchBytes_2360(matchBytes[2360]),
.io_matchBytes_2361(matchBytes[2361]),
.io_matchBytes_2362(matchBytes[2362]),
.io_matchBytes_2363(matchBytes[2363]),
.io_matchBytes_2364(matchBytes[2364]),
.io_matchBytes_2365(matchBytes[2365]),
.io_matchBytes_2366(matchBytes[2366]),
.io_matchBytes_2367(matchBytes[2367]),
.io_matchBytes_2368(matchBytes[2368]),
.io_matchBytes_2369(matchBytes[2369]),
.io_matchBytes_2370(matchBytes[2370]),
.io_matchBytes_2371(matchBytes[2371]),
.io_matchBytes_2372(matchBytes[2372]),
.io_matchBytes_2373(matchBytes[2373]),
.io_matchBytes_2374(matchBytes[2374]),
.io_matchBytes_2375(matchBytes[2375]),
.io_matchBytes_2376(matchBytes[2376]),
.io_matchBytes_2377(matchBytes[2377]),
.io_matchBytes_2378(matchBytes[2378]),
.io_matchBytes_2379(matchBytes[2379]),
.io_matchBytes_2380(matchBytes[2380]),
.io_matchBytes_2381(matchBytes[2381]),
.io_matchBytes_2382(matchBytes[2382]),
.io_matchBytes_2383(matchBytes[2383]),
.io_matchBytes_2384(matchBytes[2384]),
.io_matchBytes_2385(matchBytes[2385]),
.io_matchBytes_2386(matchBytes[2386]),
.io_matchBytes_2387(matchBytes[2387]),
.io_matchBytes_2388(matchBytes[2388]),
.io_matchBytes_2389(matchBytes[2389]),
.io_matchBytes_2390(matchBytes[2390]),
.io_matchBytes_2391(matchBytes[2391]),
.io_matchBytes_2392(matchBytes[2392]),
.io_matchBytes_2393(matchBytes[2393]),
.io_matchBytes_2394(matchBytes[2394]),
.io_matchBytes_2395(matchBytes[2395]),
.io_matchBytes_2396(matchBytes[2396]),
.io_matchBytes_2397(matchBytes[2397]),
.io_matchBytes_2398(matchBytes[2398]),
.io_matchBytes_2399(matchBytes[2399]),
.io_matchBytes_2400(matchBytes[2400]),
.io_matchBytes_2401(matchBytes[2401]),
.io_matchBytes_2402(matchBytes[2402]),
.io_matchBytes_2403(matchBytes[2403]),
.io_matchBytes_2404(matchBytes[2404]),
.io_matchBytes_2405(matchBytes[2405]),
.io_matchBytes_2406(matchBytes[2406]),
.io_matchBytes_2407(matchBytes[2407]),
.io_matchBytes_2408(matchBytes[2408]),
.io_matchBytes_2409(matchBytes[2409]),
.io_matchBytes_2410(matchBytes[2410]),
.io_matchBytes_2411(matchBytes[2411]),
.io_matchBytes_2412(matchBytes[2412]),
.io_matchBytes_2413(matchBytes[2413]),
.io_matchBytes_2414(matchBytes[2414]),
.io_matchBytes_2415(matchBytes[2415]),
.io_matchBytes_2416(matchBytes[2416]),
.io_matchBytes_2417(matchBytes[2417]),
.io_matchBytes_2418(matchBytes[2418]),
.io_matchBytes_2419(matchBytes[2419]),
.io_matchBytes_2420(matchBytes[2420]),
.io_matchBytes_2421(matchBytes[2421]),
.io_matchBytes_2422(matchBytes[2422]),
.io_matchBytes_2423(matchBytes[2423]),
.io_matchBytes_2424(matchBytes[2424]),
.io_matchBytes_2425(matchBytes[2425]),
.io_matchBytes_2426(matchBytes[2426]),
.io_matchBytes_2427(matchBytes[2427]),
.io_matchBytes_2428(matchBytes[2428]),
.io_matchBytes_2429(matchBytes[2429]),
.io_matchBytes_2430(matchBytes[2430]),
.io_matchBytes_2431(matchBytes[2431]),
.io_matchBytes_2432(matchBytes[2432]),
.io_matchBytes_2433(matchBytes[2433]),
.io_matchBytes_2434(matchBytes[2434]),
.io_matchBytes_2435(matchBytes[2435]),
.io_matchBytes_2436(matchBytes[2436]),
.io_matchBytes_2437(matchBytes[2437]),
.io_matchBytes_2438(matchBytes[2438]),
.io_matchBytes_2439(matchBytes[2439]),
.io_matchBytes_2440(matchBytes[2440]),
.io_matchBytes_2441(matchBytes[2441]),
.io_matchBytes_2442(matchBytes[2442]),
.io_matchBytes_2443(matchBytes[2443]),
.io_matchBytes_2444(matchBytes[2444]),
.io_matchBytes_2445(matchBytes[2445]),
.io_matchBytes_2446(matchBytes[2446]),
.io_matchBytes_2447(matchBytes[2447]),
.io_matchBytes_2448(matchBytes[2448]),
.io_matchBytes_2449(matchBytes[2449]),
.io_matchBytes_2450(matchBytes[2450]),
.io_matchBytes_2451(matchBytes[2451]),
.io_matchBytes_2452(matchBytes[2452]),
.io_matchBytes_2453(matchBytes[2453]),
.io_matchBytes_2454(matchBytes[2454]),
.io_matchBytes_2455(matchBytes[2455]),
.io_matchBytes_2456(matchBytes[2456]),
.io_matchBytes_2457(matchBytes[2457]),
.io_matchBytes_2458(matchBytes[2458]),
.io_matchBytes_2459(matchBytes[2459]),
.io_matchBytes_2460(matchBytes[2460]),
.io_matchBytes_2461(matchBytes[2461]),
.io_matchBytes_2462(matchBytes[2462]),
.io_matchBytes_2463(matchBytes[2463]),
.io_matchBytes_2464(matchBytes[2464]),
.io_matchBytes_2465(matchBytes[2465]),
.io_matchBytes_2466(matchBytes[2466]),
.io_matchBytes_2467(matchBytes[2467]),
.io_matchBytes_2468(matchBytes[2468]),
.io_matchBytes_2469(matchBytes[2469]),
.io_matchBytes_2470(matchBytes[2470]),
.io_matchBytes_2471(matchBytes[2471]),
.io_matchBytes_2472(matchBytes[2472]),
.io_matchBytes_2473(matchBytes[2473]),
.io_matchBytes_2474(matchBytes[2474]),
.io_matchBytes_2475(matchBytes[2475]),
.io_matchBytes_2476(matchBytes[2476]),
.io_matchBytes_2477(matchBytes[2477]),
.io_matchBytes_2478(matchBytes[2478]),
.io_matchBytes_2479(matchBytes[2479]),
.io_matchBytes_2480(matchBytes[2480]),
.io_matchBytes_2481(matchBytes[2481]),
.io_matchBytes_2482(matchBytes[2482]),
.io_matchBytes_2483(matchBytes[2483]),
.io_matchBytes_2484(matchBytes[2484]),
.io_matchBytes_2485(matchBytes[2485]),
.io_matchBytes_2486(matchBytes[2486]),
.io_matchBytes_2487(matchBytes[2487]),
.io_matchBytes_2488(matchBytes[2488]),
.io_matchBytes_2489(matchBytes[2489]),
.io_matchBytes_2490(matchBytes[2490]),
.io_matchBytes_2491(matchBytes[2491]),
.io_matchBytes_2492(matchBytes[2492]),
.io_matchBytes_2493(matchBytes[2493]),
.io_matchBytes_2494(matchBytes[2494]),
.io_matchBytes_2495(matchBytes[2495]),
.io_matchBytes_2496(matchBytes[2496]),
.io_matchBytes_2497(matchBytes[2497]),
.io_matchBytes_2498(matchBytes[2498]),
.io_matchBytes_2499(matchBytes[2499]),
.io_matchBytes_2500(matchBytes[2500]),
.io_matchBytes_2501(matchBytes[2501]),
.io_matchBytes_2502(matchBytes[2502]),
.io_matchBytes_2503(matchBytes[2503]),
.io_matchBytes_2504(matchBytes[2504]),
.io_matchBytes_2505(matchBytes[2505]),
.io_matchBytes_2506(matchBytes[2506]),
.io_matchBytes_2507(matchBytes[2507]),
.io_matchBytes_2508(matchBytes[2508]),
.io_matchBytes_2509(matchBytes[2509]),
.io_matchBytes_2510(matchBytes[2510]),
.io_matchBytes_2511(matchBytes[2511]),
.io_matchBytes_2512(matchBytes[2512]),
.io_matchBytes_2513(matchBytes[2513]),
.io_matchBytes_2514(matchBytes[2514]),
.io_matchBytes_2515(matchBytes[2515]),
.io_matchBytes_2516(matchBytes[2516]),
.io_matchBytes_2517(matchBytes[2517]),
.io_matchBytes_2518(matchBytes[2518]),
.io_matchBytes_2519(matchBytes[2519]),
.io_matchBytes_2520(matchBytes[2520]),
.io_matchBytes_2521(matchBytes[2521]),
.io_matchBytes_2522(matchBytes[2522]),
.io_matchBytes_2523(matchBytes[2523]),
.io_matchBytes_2524(matchBytes[2524]),
.io_matchBytes_2525(matchBytes[2525]),
.io_matchBytes_2526(matchBytes[2526]),
.io_matchBytes_2527(matchBytes[2527]),
.io_matchBytes_2528(matchBytes[2528]),
.io_matchBytes_2529(matchBytes[2529]),
.io_matchBytes_2530(matchBytes[2530]),
.io_matchBytes_2531(matchBytes[2531]),
.io_matchBytes_2532(matchBytes[2532]),
.io_matchBytes_2533(matchBytes[2533]),
.io_matchBytes_2534(matchBytes[2534]),
.io_matchBytes_2535(matchBytes[2535]),
.io_matchBytes_2536(matchBytes[2536]),
.io_matchBytes_2537(matchBytes[2537]),
.io_matchBytes_2538(matchBytes[2538]),
.io_matchBytes_2539(matchBytes[2539]),
.io_matchBytes_2540(matchBytes[2540]),
.io_matchBytes_2541(matchBytes[2541]),
.io_matchBytes_2542(matchBytes[2542]),
.io_matchBytes_2543(matchBytes[2543]),
.io_matchBytes_2544(matchBytes[2544]),
.io_matchBytes_2545(matchBytes[2545]),
.io_matchBytes_2546(matchBytes[2546]),
.io_matchBytes_2547(matchBytes[2547]),
.io_matchBytes_2548(matchBytes[2548]),
.io_matchBytes_2549(matchBytes[2549]),
.io_matchBytes_2550(matchBytes[2550]),
.io_matchBytes_2551(matchBytes[2551]),
.io_matchBytes_2552(matchBytes[2552]),
.io_matchBytes_2553(matchBytes[2553]),
.io_matchBytes_2554(matchBytes[2554]),
.io_matchBytes_2555(matchBytes[2555]),
.io_matchBytes_2556(matchBytes[2556]),
.io_matchBytes_2557(matchBytes[2557]),
.io_matchBytes_2558(matchBytes[2558]),
.io_matchBytes_2559(matchBytes[2559]),
.io_matchBytes_2560(matchBytes[2560]),
.io_matchBytes_2561(matchBytes[2561]),
.io_matchBytes_2562(matchBytes[2562]),
.io_matchBytes_2563(matchBytes[2563]),
.io_matchBytes_2564(matchBytes[2564]),
.io_matchBytes_2565(matchBytes[2565]),
.io_matchBytes_2566(matchBytes[2566]),
.io_matchBytes_2567(matchBytes[2567]),
.io_matchBytes_2568(matchBytes[2568]),
.io_matchBytes_2569(matchBytes[2569]),
.io_matchBytes_2570(matchBytes[2570]),
.io_matchBytes_2571(matchBytes[2571]),
.io_matchBytes_2572(matchBytes[2572]),
.io_matchBytes_2573(matchBytes[2573]),
.io_matchBytes_2574(matchBytes[2574]),
.io_matchBytes_2575(matchBytes[2575]),
.io_matchBytes_2576(matchBytes[2576]),
.io_matchBytes_2577(matchBytes[2577]),
.io_matchBytes_2578(matchBytes[2578]),
.io_matchBytes_2579(matchBytes[2579]),
.io_matchBytes_2580(matchBytes[2580]),
.io_matchBytes_2581(matchBytes[2581]),
.io_matchBytes_2582(matchBytes[2582]),
.io_matchBytes_2583(matchBytes[2583]),
.io_matchBytes_2584(matchBytes[2584]),
.io_matchBytes_2585(matchBytes[2585]),
.io_matchBytes_2586(matchBytes[2586]),
.io_matchBytes_2587(matchBytes[2587]),
.io_matchBytes_2588(matchBytes[2588]),
.io_matchBytes_2589(matchBytes[2589]),
.io_matchBytes_2590(matchBytes[2590]),
.io_matchBytes_2591(matchBytes[2591]),
.io_matchBytes_2592(matchBytes[2592]),
.io_matchBytes_2593(matchBytes[2593]),
.io_matchBytes_2594(matchBytes[2594]),
.io_matchBytes_2595(matchBytes[2595]),
.io_matchBytes_2596(matchBytes[2596]),
.io_matchBytes_2597(matchBytes[2597]),
.io_matchBytes_2598(matchBytes[2598]),
.io_matchBytes_2599(matchBytes[2599]),
.io_matchBytes_2600(matchBytes[2600]),
.io_matchBytes_2601(matchBytes[2601]),
.io_matchBytes_2602(matchBytes[2602]),
.io_matchBytes_2603(matchBytes[2603]),
.io_matchBytes_2604(matchBytes[2604]),
.io_matchBytes_2605(matchBytes[2605]),
.io_matchBytes_2606(matchBytes[2606]),
.io_matchBytes_2607(matchBytes[2607]),
.io_matchBytes_2608(matchBytes[2608]),
.io_matchBytes_2609(matchBytes[2609]),
.io_matchBytes_2610(matchBytes[2610]),
.io_matchBytes_2611(matchBytes[2611]),
.io_matchBytes_2612(matchBytes[2612]),
.io_matchBytes_2613(matchBytes[2613]),
.io_matchBytes_2614(matchBytes[2614]),
.io_matchBytes_2615(matchBytes[2615]),
.io_matchBytes_2616(matchBytes[2616]),
.io_matchBytes_2617(matchBytes[2617]),
.io_matchBytes_2618(matchBytes[2618]),
.io_matchBytes_2619(matchBytes[2619]),
.io_matchBytes_2620(matchBytes[2620]),
.io_matchBytes_2621(matchBytes[2621]),
.io_matchBytes_2622(matchBytes[2622]),
.io_matchBytes_2623(matchBytes[2623]),
.io_matchBytes_2624(matchBytes[2624]),
.io_matchBytes_2625(matchBytes[2625]),
.io_matchBytes_2626(matchBytes[2626]),
.io_matchBytes_2627(matchBytes[2627]),
.io_matchBytes_2628(matchBytes[2628]),
.io_matchBytes_2629(matchBytes[2629]),
.io_matchBytes_2630(matchBytes[2630]),
.io_matchBytes_2631(matchBytes[2631]),
.io_matchBytes_2632(matchBytes[2632]),
.io_matchBytes_2633(matchBytes[2633]),
.io_matchBytes_2634(matchBytes[2634]),
.io_matchBytes_2635(matchBytes[2635]),
.io_matchBytes_2636(matchBytes[2636]),
.io_matchBytes_2637(matchBytes[2637]),
.io_matchBytes_2638(matchBytes[2638]),
.io_matchBytes_2639(matchBytes[2639]),
.io_matchBytes_2640(matchBytes[2640]),
.io_matchBytes_2641(matchBytes[2641]),
.io_matchBytes_2642(matchBytes[2642]),
.io_matchBytes_2643(matchBytes[2643]),
.io_matchBytes_2644(matchBytes[2644]),
.io_matchBytes_2645(matchBytes[2645]),
.io_matchBytes_2646(matchBytes[2646]),
.io_matchBytes_2647(matchBytes[2647]),
.io_matchBytes_2648(matchBytes[2648]),
.io_matchBytes_2649(matchBytes[2649]),
.io_matchBytes_2650(matchBytes[2650]),
.io_matchBytes_2651(matchBytes[2651]),
.io_matchBytes_2652(matchBytes[2652]),
.io_matchBytes_2653(matchBytes[2653]),
.io_matchBytes_2654(matchBytes[2654]),
.io_matchBytes_2655(matchBytes[2655]),
.io_matchBytes_2656(matchBytes[2656]),
.io_matchBytes_2657(matchBytes[2657]),
.io_matchBytes_2658(matchBytes[2658]),
.io_matchBytes_2659(matchBytes[2659]),
.io_matchBytes_2660(matchBytes[2660]),
.io_matchBytes_2661(matchBytes[2661]),
.io_matchBytes_2662(matchBytes[2662]),
.io_matchBytes_2663(matchBytes[2663]),
.io_matchBytes_2664(matchBytes[2664]),
.io_matchBytes_2665(matchBytes[2665]),
.io_matchBytes_2666(matchBytes[2666]),
.io_matchBytes_2667(matchBytes[2667]),
.io_matchBytes_2668(matchBytes[2668]),
.io_matchBytes_2669(matchBytes[2669]),
.io_matchBytes_2670(matchBytes[2670]),
.io_matchBytes_2671(matchBytes[2671]),
.io_matchBytes_2672(matchBytes[2672]),
.io_matchBytes_2673(matchBytes[2673]),
.io_matchBytes_2674(matchBytes[2674]),
.io_matchBytes_2675(matchBytes[2675]),
.io_matchBytes_2676(matchBytes[2676]),
.io_matchBytes_2677(matchBytes[2677]),
.io_matchBytes_2678(matchBytes[2678]),
.io_matchBytes_2679(matchBytes[2679]),
.io_matchBytes_2680(matchBytes[2680]),
.io_matchBytes_2681(matchBytes[2681]),
.io_matchBytes_2682(matchBytes[2682]),
.io_matchBytes_2683(matchBytes[2683]),
.io_matchBytes_2684(matchBytes[2684]),
.io_matchBytes_2685(matchBytes[2685]),
.io_matchBytes_2686(matchBytes[2686]),
.io_matchBytes_2687(matchBytes[2687]),
.io_matchBytes_2688(matchBytes[2688]),
.io_matchBytes_2689(matchBytes[2689]),
.io_matchBytes_2690(matchBytes[2690]),
.io_matchBytes_2691(matchBytes[2691]),
.io_matchBytes_2692(matchBytes[2692]),
.io_matchBytes_2693(matchBytes[2693]),
.io_matchBytes_2694(matchBytes[2694]),
.io_matchBytes_2695(matchBytes[2695]),
.io_matchBytes_2696(matchBytes[2696]),
.io_matchBytes_2697(matchBytes[2697]),
.io_matchBytes_2698(matchBytes[2698]),
.io_matchBytes_2699(matchBytes[2699]),
.io_matchBytes_2700(matchBytes[2700]),
.io_matchBytes_2701(matchBytes[2701]),
.io_matchBytes_2702(matchBytes[2702]),
.io_matchBytes_2703(matchBytes[2703]),
.io_matchBytes_2704(matchBytes[2704]),
.io_matchBytes_2705(matchBytes[2705]),
.io_matchBytes_2706(matchBytes[2706]),
.io_matchBytes_2707(matchBytes[2707]),
.io_matchBytes_2708(matchBytes[2708]),
.io_matchBytes_2709(matchBytes[2709]),
.io_matchBytes_2710(matchBytes[2710]),
.io_matchBytes_2711(matchBytes[2711]),
.io_matchBytes_2712(matchBytes[2712]),
.io_matchBytes_2713(matchBytes[2713]),
.io_matchBytes_2714(matchBytes[2714]),
.io_matchBytes_2715(matchBytes[2715]),
.io_matchBytes_2716(matchBytes[2716]),
.io_matchBytes_2717(matchBytes[2717]),
.io_matchBytes_2718(matchBytes[2718]),
.io_matchBytes_2719(matchBytes[2719]),
.io_matchBytes_2720(matchBytes[2720]),
.io_matchBytes_2721(matchBytes[2721]),
.io_matchBytes_2722(matchBytes[2722]),
.io_matchBytes_2723(matchBytes[2723]),
.io_matchBytes_2724(matchBytes[2724]),
.io_matchBytes_2725(matchBytes[2725]),
.io_matchBytes_2726(matchBytes[2726]),
.io_matchBytes_2727(matchBytes[2727]),
.io_matchBytes_2728(matchBytes[2728]),
.io_matchBytes_2729(matchBytes[2729]),
.io_matchBytes_2730(matchBytes[2730]),
.io_matchBytes_2731(matchBytes[2731]),
.io_matchBytes_2732(matchBytes[2732]),
.io_matchBytes_2733(matchBytes[2733]),
.io_matchBytes_2734(matchBytes[2734]),
.io_matchBytes_2735(matchBytes[2735]),
.io_matchBytes_2736(matchBytes[2736]),
.io_matchBytes_2737(matchBytes[2737]),
.io_matchBytes_2738(matchBytes[2738]),
.io_matchBytes_2739(matchBytes[2739]),
.io_matchBytes_2740(matchBytes[2740]),
.io_matchBytes_2741(matchBytes[2741]),
.io_matchBytes_2742(matchBytes[2742]),
.io_matchBytes_2743(matchBytes[2743]),
.io_matchBytes_2744(matchBytes[2744]),
.io_matchBytes_2745(matchBytes[2745]),
.io_matchBytes_2746(matchBytes[2746]),
.io_matchBytes_2747(matchBytes[2747]),
.io_matchBytes_2748(matchBytes[2748]),
.io_matchBytes_2749(matchBytes[2749]),
.io_matchBytes_2750(matchBytes[2750]),
.io_matchBytes_2751(matchBytes[2751]),
.io_matchBytes_2752(matchBytes[2752]),
.io_matchBytes_2753(matchBytes[2753]),
.io_matchBytes_2754(matchBytes[2754]),
.io_matchBytes_2755(matchBytes[2755]),
.io_matchBytes_2756(matchBytes[2756]),
.io_matchBytes_2757(matchBytes[2757]),
.io_matchBytes_2758(matchBytes[2758]),
.io_matchBytes_2759(matchBytes[2759]),
.io_matchBytes_2760(matchBytes[2760]),
.io_matchBytes_2761(matchBytes[2761]),
.io_matchBytes_2762(matchBytes[2762]),
.io_matchBytes_2763(matchBytes[2763]),
.io_matchBytes_2764(matchBytes[2764]),
.io_matchBytes_2765(matchBytes[2765]),
.io_matchBytes_2766(matchBytes[2766]),
.io_matchBytes_2767(matchBytes[2767]),
.io_matchBytes_2768(matchBytes[2768]),
.io_matchBytes_2769(matchBytes[2769]),
.io_matchBytes_2770(matchBytes[2770]),
.io_matchBytes_2771(matchBytes[2771]),
.io_matchBytes_2772(matchBytes[2772]),
.io_matchBytes_2773(matchBytes[2773]),
.io_matchBytes_2774(matchBytes[2774]),
.io_matchBytes_2775(matchBytes[2775]),
.io_matchBytes_2776(matchBytes[2776]),
.io_matchBytes_2777(matchBytes[2777]),
.io_matchBytes_2778(matchBytes[2778]),
.io_matchBytes_2779(matchBytes[2779]),
.io_matchBytes_2780(matchBytes[2780]),
.io_matchBytes_2781(matchBytes[2781]),
.io_matchBytes_2782(matchBytes[2782]),
.io_matchBytes_2783(matchBytes[2783]),
.io_matchBytes_2784(matchBytes[2784]),
.io_matchBytes_2785(matchBytes[2785]),
.io_matchBytes_2786(matchBytes[2786]),
.io_matchBytes_2787(matchBytes[2787]),
.io_matchBytes_2788(matchBytes[2788]),
.io_matchBytes_2789(matchBytes[2789]),
.io_matchBytes_2790(matchBytes[2790]),
.io_matchBytes_2791(matchBytes[2791]),
.io_matchBytes_2792(matchBytes[2792]),
.io_matchBytes_2793(matchBytes[2793]),
.io_matchBytes_2794(matchBytes[2794]),
.io_matchBytes_2795(matchBytes[2795]),
.io_matchBytes_2796(matchBytes[2796]),
.io_matchBytes_2797(matchBytes[2797]),
.io_matchBytes_2798(matchBytes[2798]),
.io_matchBytes_2799(matchBytes[2799]),
.io_matchBytes_2800(matchBytes[2800]),
.io_matchBytes_2801(matchBytes[2801]),
.io_matchBytes_2802(matchBytes[2802]),
.io_matchBytes_2803(matchBytes[2803]),
.io_matchBytes_2804(matchBytes[2804]),
.io_matchBytes_2805(matchBytes[2805]),
.io_matchBytes_2806(matchBytes[2806]),
.io_matchBytes_2807(matchBytes[2807]),
.io_matchBytes_2808(matchBytes[2808]),
.io_matchBytes_2809(matchBytes[2809]),
.io_matchBytes_2810(matchBytes[2810]),
.io_matchBytes_2811(matchBytes[2811]),
.io_matchBytes_2812(matchBytes[2812]),
.io_matchBytes_2813(matchBytes[2813]),
.io_matchBytes_2814(matchBytes[2814]),
.io_matchBytes_2815(matchBytes[2815]),
.io_matchBytes_2816(matchBytes[2816]),
.io_matchBytes_2817(matchBytes[2817]),
.io_matchBytes_2818(matchBytes[2818]),
.io_matchBytes_2819(matchBytes[2819]),
.io_matchBytes_2820(matchBytes[2820]),
.io_matchBytes_2821(matchBytes[2821]),
.io_matchBytes_2822(matchBytes[2822]),
.io_matchBytes_2823(matchBytes[2823]),
.io_matchBytes_2824(matchBytes[2824]),
.io_matchBytes_2825(matchBytes[2825]),
.io_matchBytes_2826(matchBytes[2826]),
.io_matchBytes_2827(matchBytes[2827]),
.io_matchBytes_2828(matchBytes[2828]),
.io_matchBytes_2829(matchBytes[2829]),
.io_matchBytes_2830(matchBytes[2830]),
.io_matchBytes_2831(matchBytes[2831]),
.io_matchBytes_2832(matchBytes[2832]),
.io_matchBytes_2833(matchBytes[2833]),
.io_matchBytes_2834(matchBytes[2834]),
.io_matchBytes_2835(matchBytes[2835]),
.io_matchBytes_2836(matchBytes[2836]),
.io_matchBytes_2837(matchBytes[2837]),
.io_matchBytes_2838(matchBytes[2838]),
.io_matchBytes_2839(matchBytes[2839]),
.io_matchBytes_2840(matchBytes[2840]),
.io_matchBytes_2841(matchBytes[2841]),
.io_matchBytes_2842(matchBytes[2842]),
.io_matchBytes_2843(matchBytes[2843]),
.io_matchBytes_2844(matchBytes[2844]),
.io_matchBytes_2845(matchBytes[2845]),
.io_matchBytes_2846(matchBytes[2846]),
.io_matchBytes_2847(matchBytes[2847]),
.io_matchBytes_2848(matchBytes[2848]),
.io_matchBytes_2849(matchBytes[2849]),
.io_matchBytes_2850(matchBytes[2850]),
.io_matchBytes_2851(matchBytes[2851]),
.io_matchBytes_2852(matchBytes[2852]),
.io_matchBytes_2853(matchBytes[2853]),
.io_matchBytes_2854(matchBytes[2854]),
.io_matchBytes_2855(matchBytes[2855]),
.io_matchBytes_2856(matchBytes[2856]),
.io_matchBytes_2857(matchBytes[2857]),
.io_matchBytes_2858(matchBytes[2858]),
.io_matchBytes_2859(matchBytes[2859]),
.io_matchBytes_2860(matchBytes[2860]),
.io_matchBytes_2861(matchBytes[2861]),
.io_matchBytes_2862(matchBytes[2862]),
.io_matchBytes_2863(matchBytes[2863]),
.io_matchBytes_2864(matchBytes[2864]),
.io_matchBytes_2865(matchBytes[2865]),
.io_matchBytes_2866(matchBytes[2866]),
.io_matchBytes_2867(matchBytes[2867]),
.io_matchBytes_2868(matchBytes[2868]),
.io_matchBytes_2869(matchBytes[2869]),
.io_matchBytes_2870(matchBytes[2870]),
.io_matchBytes_2871(matchBytes[2871]),
.io_matchBytes_2872(matchBytes[2872]),
.io_matchBytes_2873(matchBytes[2873]),
.io_matchBytes_2874(matchBytes[2874]),
.io_matchBytes_2875(matchBytes[2875]),
.io_matchBytes_2876(matchBytes[2876]),
.io_matchBytes_2877(matchBytes[2877]),
.io_matchBytes_2878(matchBytes[2878]),
.io_matchBytes_2879(matchBytes[2879]),
.io_matchBytes_2880(matchBytes[2880]),
.io_matchBytes_2881(matchBytes[2881]),
.io_matchBytes_2882(matchBytes[2882]),
.io_matchBytes_2883(matchBytes[2883]),
.io_matchBytes_2884(matchBytes[2884]),
.io_matchBytes_2885(matchBytes[2885]),
.io_matchBytes_2886(matchBytes[2886]),
.io_matchBytes_2887(matchBytes[2887]),
.io_matchBytes_2888(matchBytes[2888]),
.io_matchBytes_2889(matchBytes[2889]),
.io_matchBytes_2890(matchBytes[2890]),
.io_matchBytes_2891(matchBytes[2891]),
.io_matchBytes_2892(matchBytes[2892]),
.io_matchBytes_2893(matchBytes[2893]),
.io_matchBytes_2894(matchBytes[2894]),
.io_matchBytes_2895(matchBytes[2895]),
.io_matchBytes_2896(matchBytes[2896]),
.io_matchBytes_2897(matchBytes[2897]),
.io_matchBytes_2898(matchBytes[2898]),
.io_matchBytes_2899(matchBytes[2899]),
.io_matchBytes_2900(matchBytes[2900]),
.io_matchBytes_2901(matchBytes[2901]),
.io_matchBytes_2902(matchBytes[2902]),
.io_matchBytes_2903(matchBytes[2903]),
.io_matchBytes_2904(matchBytes[2904]),
.io_matchBytes_2905(matchBytes[2905]),
.io_matchBytes_2906(matchBytes[2906]),
.io_matchBytes_2907(matchBytes[2907]),
.io_matchBytes_2908(matchBytes[2908]),
.io_matchBytes_2909(matchBytes[2909]),
.io_matchBytes_2910(matchBytes[2910]),
.io_matchBytes_2911(matchBytes[2911]),
.io_matchBytes_2912(matchBytes[2912]),
.io_matchBytes_2913(matchBytes[2913]),
.io_matchBytes_2914(matchBytes[2914]),
.io_matchBytes_2915(matchBytes[2915]),
.io_matchBytes_2916(matchBytes[2916]),
.io_matchBytes_2917(matchBytes[2917]),
.io_matchBytes_2918(matchBytes[2918]),
.io_matchBytes_2919(matchBytes[2919]),
.io_matchBytes_2920(matchBytes[2920]),
.io_matchBytes_2921(matchBytes[2921]),
.io_matchBytes_2922(matchBytes[2922]),
.io_matchBytes_2923(matchBytes[2923]),
.io_matchBytes_2924(matchBytes[2924]),
.io_matchBytes_2925(matchBytes[2925]),
.io_matchBytes_2926(matchBytes[2926]),
.io_matchBytes_2927(matchBytes[2927]),
.io_matchBytes_2928(matchBytes[2928]),
.io_matchBytes_2929(matchBytes[2929]),
.io_matchBytes_2930(matchBytes[2930]),
.io_matchBytes_2931(matchBytes[2931]),
.io_matchBytes_2932(matchBytes[2932]),
.io_matchBytes_2933(matchBytes[2933]),
.io_matchBytes_2934(matchBytes[2934]),
.io_matchBytes_2935(matchBytes[2935]),
.io_matchBytes_2936(matchBytes[2936]),
.io_matchBytes_2937(matchBytes[2937]),
.io_matchBytes_2938(matchBytes[2938]),
.io_matchBytes_2939(matchBytes[2939]),
.io_matchBytes_2940(matchBytes[2940]),
.io_matchBytes_2941(matchBytes[2941]),
.io_matchBytes_2942(matchBytes[2942]),
.io_matchBytes_2943(matchBytes[2943]),
.io_matchBytes_2944(matchBytes[2944]),
.io_matchBytes_2945(matchBytes[2945]),
.io_matchBytes_2946(matchBytes[2946]),
.io_matchBytes_2947(matchBytes[2947]),
.io_matchBytes_2948(matchBytes[2948]),
.io_matchBytes_2949(matchBytes[2949]),
.io_matchBytes_2950(matchBytes[2950]),
.io_matchBytes_2951(matchBytes[2951]),
.io_matchBytes_2952(matchBytes[2952]),
.io_matchBytes_2953(matchBytes[2953]),
.io_matchBytes_2954(matchBytes[2954]),
.io_matchBytes_2955(matchBytes[2955]),
.io_matchBytes_2956(matchBytes[2956]),
.io_matchBytes_2957(matchBytes[2957]),
.io_matchBytes_2958(matchBytes[2958]),
.io_matchBytes_2959(matchBytes[2959]),
.io_matchBytes_2960(matchBytes[2960]),
.io_matchBytes_2961(matchBytes[2961]),
.io_matchBytes_2962(matchBytes[2962]),
.io_matchBytes_2963(matchBytes[2963]),
.io_matchBytes_2964(matchBytes[2964]),
.io_matchBytes_2965(matchBytes[2965]),
.io_matchBytes_2966(matchBytes[2966]),
.io_matchBytes_2967(matchBytes[2967]),
.io_matchBytes_2968(matchBytes[2968]),
.io_matchBytes_2969(matchBytes[2969]),
.io_matchBytes_2970(matchBytes[2970]),
.io_matchBytes_2971(matchBytes[2971]),
.io_matchBytes_2972(matchBytes[2972]),
.io_matchBytes_2973(matchBytes[2973]),
.io_matchBytes_2974(matchBytes[2974]),
.io_matchBytes_2975(matchBytes[2975]),
.io_matchBytes_2976(matchBytes[2976]),
.io_matchBytes_2977(matchBytes[2977]),
.io_matchBytes_2978(matchBytes[2978]),
.io_matchBytes_2979(matchBytes[2979]),
.io_matchBytes_2980(matchBytes[2980]),
.io_matchBytes_2981(matchBytes[2981]),
.io_matchBytes_2982(matchBytes[2982]),
.io_matchBytes_2983(matchBytes[2983]),
.io_matchBytes_2984(matchBytes[2984]),
.io_matchBytes_2985(matchBytes[2985]),
.io_matchBytes_2986(matchBytes[2986]),
.io_matchBytes_2987(matchBytes[2987]),
.io_matchBytes_2988(matchBytes[2988]),
.io_matchBytes_2989(matchBytes[2989]),
.io_matchBytes_2990(matchBytes[2990]),
.io_matchBytes_2991(matchBytes[2991]),
.io_matchBytes_2992(matchBytes[2992]),
.io_matchBytes_2993(matchBytes[2993]),
.io_matchBytes_2994(matchBytes[2994]),
.io_matchBytes_2995(matchBytes[2995]),
.io_matchBytes_2996(matchBytes[2996]),
.io_matchBytes_2997(matchBytes[2997]),
.io_matchBytes_2998(matchBytes[2998]),
.io_matchBytes_2999(matchBytes[2999]),
.io_matchBytes_3000(matchBytes[3000]),
.io_matchBytes_3001(matchBytes[3001]),
.io_matchBytes_3002(matchBytes[3002]),
.io_matchBytes_3003(matchBytes[3003]),
.io_matchBytes_3004(matchBytes[3004]),
.io_matchBytes_3005(matchBytes[3005]),
.io_matchBytes_3006(matchBytes[3006]),
.io_matchBytes_3007(matchBytes[3007]),
.io_matchBytes_3008(matchBytes[3008]),
.io_matchBytes_3009(matchBytes[3009]),
.io_matchBytes_3010(matchBytes[3010]),
.io_matchBytes_3011(matchBytes[3011]),
.io_matchBytes_3012(matchBytes[3012]),
.io_matchBytes_3013(matchBytes[3013]),
.io_matchBytes_3014(matchBytes[3014]),
.io_matchBytes_3015(matchBytes[3015]),
.io_matchBytes_3016(matchBytes[3016]),
.io_matchBytes_3017(matchBytes[3017]),
.io_matchBytes_3018(matchBytes[3018]),
.io_matchBytes_3019(matchBytes[3019]),
.io_matchBytes_3020(matchBytes[3020]),
.io_matchBytes_3021(matchBytes[3021]),
.io_matchBytes_3022(matchBytes[3022]),
.io_matchBytes_3023(matchBytes[3023]),
.io_matchBytes_3024(matchBytes[3024]),
.io_matchBytes_3025(matchBytes[3025]),
.io_matchBytes_3026(matchBytes[3026]),
.io_matchBytes_3027(matchBytes[3027]),
.io_matchBytes_3028(matchBytes[3028]),
.io_matchBytes_3029(matchBytes[3029]),
.io_matchBytes_3030(matchBytes[3030]),
.io_matchBytes_3031(matchBytes[3031]),
.io_matchBytes_3032(matchBytes[3032]),
.io_matchBytes_3033(matchBytes[3033]),
.io_matchBytes_3034(matchBytes[3034]),
.io_matchBytes_3035(matchBytes[3035]),
.io_matchBytes_3036(matchBytes[3036]),
.io_matchBytes_3037(matchBytes[3037]),
.io_matchBytes_3038(matchBytes[3038]),
.io_matchBytes_3039(matchBytes[3039]),
.io_matchBytes_3040(matchBytes[3040]),
.io_matchBytes_3041(matchBytes[3041]),
.io_matchBytes_3042(matchBytes[3042]),
.io_matchBytes_3043(matchBytes[3043]),
.io_matchBytes_3044(matchBytes[3044]),
.io_matchBytes_3045(matchBytes[3045]),
.io_matchBytes_3046(matchBytes[3046]),
.io_matchBytes_3047(matchBytes[3047]),
.io_matchBytes_3048(matchBytes[3048]),
.io_matchBytes_3049(matchBytes[3049]),
.io_matchBytes_3050(matchBytes[3050]),
.io_matchBytes_3051(matchBytes[3051]),
.io_matchBytes_3052(matchBytes[3052]),
.io_matchBytes_3053(matchBytes[3053]),
.io_matchBytes_3054(matchBytes[3054]),
.io_matchBytes_3055(matchBytes[3055]),
.io_matchBytes_3056(matchBytes[3056]),
.io_matchBytes_3057(matchBytes[3057]),
.io_matchBytes_3058(matchBytes[3058]),
.io_matchBytes_3059(matchBytes[3059]),
.io_matchBytes_3060(matchBytes[3060]),
.io_matchBytes_3061(matchBytes[3061]),
.io_matchBytes_3062(matchBytes[3062]),
.io_matchBytes_3063(matchBytes[3063]),
.io_matchBytes_3064(matchBytes[3064]),
.io_matchBytes_3065(matchBytes[3065]),
.io_matchBytes_3066(matchBytes[3066]),
.io_matchBytes_3067(matchBytes[3067]),
.io_matchBytes_3068(matchBytes[3068]),
.io_matchBytes_3069(matchBytes[3069]),
.io_matchBytes_3070(matchBytes[3070]),
.io_matchBytes_3071(matchBytes[3071]),
.io_matchBytes_3072(matchBytes[3072]),
.io_matchBytes_3073(matchBytes[3073]),
.io_matchBytes_3074(matchBytes[3074]),
.io_matchBytes_3075(matchBytes[3075]),
.io_matchBytes_3076(matchBytes[3076]),
.io_matchBytes_3077(matchBytes[3077]),
.io_matchBytes_3078(matchBytes[3078]),
.io_matchBytes_3079(matchBytes[3079]),
.io_matchBytes_3080(matchBytes[3080]),
.io_matchBytes_3081(matchBytes[3081]),
.io_matchBytes_3082(matchBytes[3082]),
.io_matchBytes_3083(matchBytes[3083]),
.io_matchBytes_3084(matchBytes[3084]),
.io_matchBytes_3085(matchBytes[3085]),
.io_matchBytes_3086(matchBytes[3086]),
.io_matchBytes_3087(matchBytes[3087]),
.io_matchBytes_3088(matchBytes[3088]),
.io_matchBytes_3089(matchBytes[3089]),
.io_matchBytes_3090(matchBytes[3090]),
.io_matchBytes_3091(matchBytes[3091]),
.io_matchBytes_3092(matchBytes[3092]),
.io_matchBytes_3093(matchBytes[3093]),
.io_matchBytes_3094(matchBytes[3094]),
.io_matchBytes_3095(matchBytes[3095]),
.io_matchBytes_3096(matchBytes[3096]),
.io_matchBytes_3097(matchBytes[3097]),
.io_matchBytes_3098(matchBytes[3098]),
.io_matchBytes_3099(matchBytes[3099]),
.io_matchBytes_3100(matchBytes[3100]),
.io_matchBytes_3101(matchBytes[3101]),
.io_matchBytes_3102(matchBytes[3102]),
.io_matchBytes_3103(matchBytes[3103]),
.io_matchBytes_3104(matchBytes[3104]),
.io_matchBytes_3105(matchBytes[3105]),
.io_matchBytes_3106(matchBytes[3106]),
.io_matchBytes_3107(matchBytes[3107]),
.io_matchBytes_3108(matchBytes[3108]),
.io_matchBytes_3109(matchBytes[3109]),
.io_matchBytes_3110(matchBytes[3110]),
.io_matchBytes_3111(matchBytes[3111]),
.io_matchBytes_3112(matchBytes[3112]),
.io_matchBytes_3113(matchBytes[3113]),
.io_matchBytes_3114(matchBytes[3114]),
.io_matchBytes_3115(matchBytes[3115]),
.io_matchBytes_3116(matchBytes[3116]),
.io_matchBytes_3117(matchBytes[3117]),
.io_matchBytes_3118(matchBytes[3118]),
.io_matchBytes_3119(matchBytes[3119]),
.io_matchBytes_3120(matchBytes[3120]),
.io_matchBytes_3121(matchBytes[3121]),
.io_matchBytes_3122(matchBytes[3122]),
.io_matchBytes_3123(matchBytes[3123]),
.io_matchBytes_3124(matchBytes[3124]),
.io_matchBytes_3125(matchBytes[3125]),
.io_matchBytes_3126(matchBytes[3126]),
.io_matchBytes_3127(matchBytes[3127]),
.io_matchBytes_3128(matchBytes[3128]),
.io_matchBytes_3129(matchBytes[3129]),
.io_matchBytes_3130(matchBytes[3130]),
.io_matchBytes_3131(matchBytes[3131]),
.io_matchBytes_3132(matchBytes[3132]),
.io_matchBytes_3133(matchBytes[3133]),
.io_matchBytes_3134(matchBytes[3134]),
.io_matchBytes_3135(matchBytes[3135]),
.io_matchBytes_3136(matchBytes[3136]),
.io_matchBytes_3137(matchBytes[3137]),
.io_matchBytes_3138(matchBytes[3138]),
.io_matchBytes_3139(matchBytes[3139]),
.io_matchBytes_3140(matchBytes[3140]),
.io_matchBytes_3141(matchBytes[3141]),
.io_matchBytes_3142(matchBytes[3142]),
.io_matchBytes_3143(matchBytes[3143]),
.io_matchBytes_3144(matchBytes[3144]),
.io_matchBytes_3145(matchBytes[3145]),
.io_matchBytes_3146(matchBytes[3146]),
.io_matchBytes_3147(matchBytes[3147]),
.io_matchBytes_3148(matchBytes[3148]),
.io_matchBytes_3149(matchBytes[3149]),
.io_matchBytes_3150(matchBytes[3150]),
.io_matchBytes_3151(matchBytes[3151]),
.io_matchBytes_3152(matchBytes[3152]),
.io_matchBytes_3153(matchBytes[3153]),
.io_matchBytes_3154(matchBytes[3154]),
.io_matchBytes_3155(matchBytes[3155]),
.io_matchBytes_3156(matchBytes[3156]),
.io_matchBytes_3157(matchBytes[3157]),
.io_matchBytes_3158(matchBytes[3158]),
.io_matchBytes_3159(matchBytes[3159]),
.io_matchBytes_3160(matchBytes[3160]),
.io_matchBytes_3161(matchBytes[3161]),
.io_matchBytes_3162(matchBytes[3162]),
.io_matchBytes_3163(matchBytes[3163]),
.io_matchBytes_3164(matchBytes[3164]),
.io_matchBytes_3165(matchBytes[3165]),
.io_matchBytes_3166(matchBytes[3166]),
.io_matchBytes_3167(matchBytes[3167]),
.io_matchBytes_3168(matchBytes[3168]),
.io_matchBytes_3169(matchBytes[3169]),
.io_matchBytes_3170(matchBytes[3170]),
.io_matchBytes_3171(matchBytes[3171]),
.io_matchBytes_3172(matchBytes[3172]),
.io_matchBytes_3173(matchBytes[3173]),
.io_matchBytes_3174(matchBytes[3174]),
.io_matchBytes_3175(matchBytes[3175]),
.io_matchBytes_3176(matchBytes[3176]),
.io_matchBytes_3177(matchBytes[3177]),
.io_matchBytes_3178(matchBytes[3178]),
.io_matchBytes_3179(matchBytes[3179]),
.io_matchBytes_3180(matchBytes[3180]),
.io_matchBytes_3181(matchBytes[3181]),
.io_matchBytes_3182(matchBytes[3182]),
.io_matchBytes_3183(matchBytes[3183]),
.io_matchBytes_3184(matchBytes[3184]),
.io_matchBytes_3185(matchBytes[3185]),
.io_matchBytes_3186(matchBytes[3186]),
.io_matchBytes_3187(matchBytes[3187]),
.io_matchBytes_3188(matchBytes[3188]),
.io_matchBytes_3189(matchBytes[3189]),
.io_matchBytes_3190(matchBytes[3190]),
.io_matchBytes_3191(matchBytes[3191]),
.io_matchBytes_3192(matchBytes[3192]),
.io_matchBytes_3193(matchBytes[3193]),
.io_matchBytes_3194(matchBytes[3194]),
.io_matchBytes_3195(matchBytes[3195]),
.io_matchBytes_3196(matchBytes[3196]),
.io_matchBytes_3197(matchBytes[3197]),
.io_matchBytes_3198(matchBytes[3198]),
.io_matchBytes_3199(matchBytes[3199]),
.io_matchBytes_3200(matchBytes[3200]),
.io_matchBytes_3201(matchBytes[3201]),
.io_matchBytes_3202(matchBytes[3202]),
.io_matchBytes_3203(matchBytes[3203]),
.io_matchBytes_3204(matchBytes[3204]),
.io_matchBytes_3205(matchBytes[3205]),
.io_matchBytes_3206(matchBytes[3206]),
.io_matchBytes_3207(matchBytes[3207]),
.io_matchBytes_3208(matchBytes[3208]),
.io_matchBytes_3209(matchBytes[3209]),
.io_matchBytes_3210(matchBytes[3210]),
.io_matchBytes_3211(matchBytes[3211]),
.io_matchBytes_3212(matchBytes[3212]),
.io_matchBytes_3213(matchBytes[3213]),
.io_matchBytes_3214(matchBytes[3214]),
.io_matchBytes_3215(matchBytes[3215]),
.io_matchBytes_3216(matchBytes[3216]),
.io_matchBytes_3217(matchBytes[3217]),
.io_matchBytes_3218(matchBytes[3218]),
.io_matchBytes_3219(matchBytes[3219]),
.io_matchBytes_3220(matchBytes[3220]),
.io_matchBytes_3221(matchBytes[3221]),
.io_matchBytes_3222(matchBytes[3222]),
.io_matchBytes_3223(matchBytes[3223]),
.io_matchBytes_3224(matchBytes[3224]),
.io_matchBytes_3225(matchBytes[3225]),
.io_matchBytes_3226(matchBytes[3226]),
.io_matchBytes_3227(matchBytes[3227]),
.io_matchBytes_3228(matchBytes[3228]),
.io_matchBytes_3229(matchBytes[3229]),
.io_matchBytes_3230(matchBytes[3230]),
.io_matchBytes_3231(matchBytes[3231]),
.io_matchBytes_3232(matchBytes[3232]),
.io_matchBytes_3233(matchBytes[3233]),
.io_matchBytes_3234(matchBytes[3234]),
.io_matchBytes_3235(matchBytes[3235]),
.io_matchBytes_3236(matchBytes[3236]),
.io_matchBytes_3237(matchBytes[3237]),
.io_matchBytes_3238(matchBytes[3238]),
.io_matchBytes_3239(matchBytes[3239]),
.io_matchBytes_3240(matchBytes[3240]),
.io_matchBytes_3241(matchBytes[3241]),
.io_matchBytes_3242(matchBytes[3242]),
.io_matchBytes_3243(matchBytes[3243]),
.io_matchBytes_3244(matchBytes[3244]),
.io_matchBytes_3245(matchBytes[3245]),
.io_matchBytes_3246(matchBytes[3246]),
.io_matchBytes_3247(matchBytes[3247]),
.io_matchBytes_3248(matchBytes[3248]),
.io_matchBytes_3249(matchBytes[3249]),
.io_matchBytes_3250(matchBytes[3250]),
.io_matchBytes_3251(matchBytes[3251]),
.io_matchBytes_3252(matchBytes[3252]),
.io_matchBytes_3253(matchBytes[3253]),
.io_matchBytes_3254(matchBytes[3254]),
.io_matchBytes_3255(matchBytes[3255]),
.io_matchBytes_3256(matchBytes[3256]),
.io_matchBytes_3257(matchBytes[3257]),
.io_matchBytes_3258(matchBytes[3258]),
.io_matchBytes_3259(matchBytes[3259]),
.io_matchBytes_3260(matchBytes[3260]),
.io_matchBytes_3261(matchBytes[3261]),
.io_matchBytes_3262(matchBytes[3262]),
.io_matchBytes_3263(matchBytes[3263]),
.io_matchBytes_3264(matchBytes[3264]),
.io_matchBytes_3265(matchBytes[3265]),
.io_matchBytes_3266(matchBytes[3266]),
.io_matchBytes_3267(matchBytes[3267]),
.io_matchBytes_3268(matchBytes[3268]),
.io_matchBytes_3269(matchBytes[3269]),
.io_matchBytes_3270(matchBytes[3270]),
.io_matchBytes_3271(matchBytes[3271]),
.io_matchBytes_3272(matchBytes[3272]),
.io_matchBytes_3273(matchBytes[3273]),
.io_matchBytes_3274(matchBytes[3274]),
.io_matchBytes_3275(matchBytes[3275]),
.io_matchBytes_3276(matchBytes[3276]),
.io_matchBytes_3277(matchBytes[3277]),
.io_matchBytes_3278(matchBytes[3278]),
.io_matchBytes_3279(matchBytes[3279]),
.io_matchBytes_3280(matchBytes[3280]),
.io_matchBytes_3281(matchBytes[3281]),
.io_matchBytes_3282(matchBytes[3282]),
.io_matchBytes_3283(matchBytes[3283]),
.io_matchBytes_3284(matchBytes[3284]),
.io_matchBytes_3285(matchBytes[3285]),
.io_matchBytes_3286(matchBytes[3286]),
.io_matchBytes_3287(matchBytes[3287]),
.io_matchBytes_3288(matchBytes[3288]),
.io_matchBytes_3289(matchBytes[3289]),
.io_matchBytes_3290(matchBytes[3290]),
.io_matchBytes_3291(matchBytes[3291]),
.io_matchBytes_3292(matchBytes[3292]),
.io_matchBytes_3293(matchBytes[3293]),
.io_matchBytes_3294(matchBytes[3294]),
.io_matchBytes_3295(matchBytes[3295]),
.io_matchBytes_3296(matchBytes[3296]),
.io_matchBytes_3297(matchBytes[3297]),
.io_matchBytes_3298(matchBytes[3298]),
.io_matchBytes_3299(matchBytes[3299]),
.io_matchBytes_3300(matchBytes[3300]),
.io_matchBytes_3301(matchBytes[3301]),
.io_matchBytes_3302(matchBytes[3302]),
.io_matchBytes_3303(matchBytes[3303]),
.io_matchBytes_3304(matchBytes[3304]),
.io_matchBytes_3305(matchBytes[3305]),
.io_matchBytes_3306(matchBytes[3306]),
.io_matchBytes_3307(matchBytes[3307]),
.io_matchBytes_3308(matchBytes[3308]),
.io_matchBytes_3309(matchBytes[3309]),
.io_matchBytes_3310(matchBytes[3310]),
.io_matchBytes_3311(matchBytes[3311]),
.io_matchBytes_3312(matchBytes[3312]),
.io_matchBytes_3313(matchBytes[3313]),
.io_matchBytes_3314(matchBytes[3314]),
.io_matchBytes_3315(matchBytes[3315]),
.io_matchBytes_3316(matchBytes[3316]),
.io_matchBytes_3317(matchBytes[3317]),
.io_matchBytes_3318(matchBytes[3318]),
.io_matchBytes_3319(matchBytes[3319]),
.io_matchBytes_3320(matchBytes[3320]),
.io_matchBytes_3321(matchBytes[3321]),
.io_matchBytes_3322(matchBytes[3322]),
.io_matchBytes_3323(matchBytes[3323]),
.io_matchBytes_3324(matchBytes[3324]),
.io_matchBytes_3325(matchBytes[3325]),
.io_matchBytes_3326(matchBytes[3326]),
.io_matchBytes_3327(matchBytes[3327]),
.io_matchBytes_3328(matchBytes[3328]),
.io_matchBytes_3329(matchBytes[3329]),
.io_matchBytes_3330(matchBytes[3330]),
.io_matchBytes_3331(matchBytes[3331]),
.io_matchBytes_3332(matchBytes[3332]),
.io_matchBytes_3333(matchBytes[3333]),
.io_matchBytes_3334(matchBytes[3334]),
.io_matchBytes_3335(matchBytes[3335]),
.io_matchBytes_3336(matchBytes[3336]),
.io_matchBytes_3337(matchBytes[3337]),
.io_matchBytes_3338(matchBytes[3338]),
.io_matchBytes_3339(matchBytes[3339]),
.io_matchBytes_3340(matchBytes[3340]),
.io_matchBytes_3341(matchBytes[3341]),
.io_matchBytes_3342(matchBytes[3342]),
.io_matchBytes_3343(matchBytes[3343]),
.io_matchBytes_3344(matchBytes[3344]),
.io_matchBytes_3345(matchBytes[3345]),
.io_matchBytes_3346(matchBytes[3346]),
.io_matchBytes_3347(matchBytes[3347]),
.io_matchBytes_3348(matchBytes[3348]),
.io_matchBytes_3349(matchBytes[3349]),
.io_matchBytes_3350(matchBytes[3350]),
.io_matchBytes_3351(matchBytes[3351]),
.io_matchBytes_3352(matchBytes[3352]),
.io_matchBytes_3353(matchBytes[3353]),
.io_matchBytes_3354(matchBytes[3354]),
.io_matchBytes_3355(matchBytes[3355]),
.io_matchBytes_3356(matchBytes[3356]),
.io_matchBytes_3357(matchBytes[3357]),
.io_matchBytes_3358(matchBytes[3358]),
.io_matchBytes_3359(matchBytes[3359]),
.io_matchBytes_3360(matchBytes[3360]),
.io_matchBytes_3361(matchBytes[3361]),
.io_matchBytes_3362(matchBytes[3362]),
.io_matchBytes_3363(matchBytes[3363]),
.io_matchBytes_3364(matchBytes[3364]),
.io_matchBytes_3365(matchBytes[3365]),
.io_matchBytes_3366(matchBytes[3366]),
.io_matchBytes_3367(matchBytes[3367]),
.io_matchBytes_3368(matchBytes[3368]),
.io_matchBytes_3369(matchBytes[3369]),
.io_matchBytes_3370(matchBytes[3370]),
.io_matchBytes_3371(matchBytes[3371]),
.io_matchBytes_3372(matchBytes[3372]),
.io_matchBytes_3373(matchBytes[3373]),
.io_matchBytes_3374(matchBytes[3374]),
.io_matchBytes_3375(matchBytes[3375]),
.io_matchBytes_3376(matchBytes[3376]),
.io_matchBytes_3377(matchBytes[3377]),
.io_matchBytes_3378(matchBytes[3378]),
.io_matchBytes_3379(matchBytes[3379]),
.io_matchBytes_3380(matchBytes[3380]),
.io_matchBytes_3381(matchBytes[3381]),
.io_matchBytes_3382(matchBytes[3382]),
.io_matchBytes_3383(matchBytes[3383]),
.io_matchBytes_3384(matchBytes[3384]),
.io_matchBytes_3385(matchBytes[3385]),
.io_matchBytes_3386(matchBytes[3386]),
.io_matchBytes_3387(matchBytes[3387]),
.io_matchBytes_3388(matchBytes[3388]),
.io_matchBytes_3389(matchBytes[3389]),
.io_matchBytes_3390(matchBytes[3390]),
.io_matchBytes_3391(matchBytes[3391]),
.io_matchBytes_3392(matchBytes[3392]),
.io_matchBytes_3393(matchBytes[3393]),
.io_matchBytes_3394(matchBytes[3394]),
.io_matchBytes_3395(matchBytes[3395]),
.io_matchBytes_3396(matchBytes[3396]),
.io_matchBytes_3397(matchBytes[3397]),
.io_matchBytes_3398(matchBytes[3398]),
.io_matchBytes_3399(matchBytes[3399]),
.io_matchBytes_3400(matchBytes[3400]),
.io_matchBytes_3401(matchBytes[3401]),
.io_matchBytes_3402(matchBytes[3402]),
.io_matchBytes_3403(matchBytes[3403]),
.io_matchBytes_3404(matchBytes[3404]),
.io_matchBytes_3405(matchBytes[3405]),
.io_matchBytes_3406(matchBytes[3406]),
.io_matchBytes_3407(matchBytes[3407]),
.io_matchBytes_3408(matchBytes[3408]),
.io_matchBytes_3409(matchBytes[3409]),
.io_matchBytes_3410(matchBytes[3410]),
.io_matchBytes_3411(matchBytes[3411]),
.io_matchBytes_3412(matchBytes[3412]),
.io_matchBytes_3413(matchBytes[3413]),
.io_matchBytes_3414(matchBytes[3414]),
.io_matchBytes_3415(matchBytes[3415]),
.io_matchBytes_3416(matchBytes[3416]),
.io_matchBytes_3417(matchBytes[3417]),
.io_matchBytes_3418(matchBytes[3418]),
.io_matchBytes_3419(matchBytes[3419]),
.io_matchBytes_3420(matchBytes[3420]),
.io_matchBytes_3421(matchBytes[3421]),
.io_matchBytes_3422(matchBytes[3422]),
.io_matchBytes_3423(matchBytes[3423]),
.io_matchBytes_3424(matchBytes[3424]),
.io_matchBytes_3425(matchBytes[3425]),
.io_matchBytes_3426(matchBytes[3426]),
.io_matchBytes_3427(matchBytes[3427]),
.io_matchBytes_3428(matchBytes[3428]),
.io_matchBytes_3429(matchBytes[3429]),
.io_matchBytes_3430(matchBytes[3430]),
.io_matchBytes_3431(matchBytes[3431]),
.io_matchBytes_3432(matchBytes[3432]),
.io_matchBytes_3433(matchBytes[3433]),
.io_matchBytes_3434(matchBytes[3434]),
.io_matchBytes_3435(matchBytes[3435]),
.io_matchBytes_3436(matchBytes[3436]),
.io_matchBytes_3437(matchBytes[3437]),
.io_matchBytes_3438(matchBytes[3438]),
.io_matchBytes_3439(matchBytes[3439]),
.io_matchBytes_3440(matchBytes[3440]),
.io_matchBytes_3441(matchBytes[3441]),
.io_matchBytes_3442(matchBytes[3442]),
.io_matchBytes_3443(matchBytes[3443]),
.io_matchBytes_3444(matchBytes[3444]),
.io_matchBytes_3445(matchBytes[3445]),
.io_matchBytes_3446(matchBytes[3446]),
.io_matchBytes_3447(matchBytes[3447]),
.io_matchBytes_3448(matchBytes[3448]),
.io_matchBytes_3449(matchBytes[3449]),
.io_matchBytes_3450(matchBytes[3450]),
.io_matchBytes_3451(matchBytes[3451]),
.io_matchBytes_3452(matchBytes[3452]),
.io_matchBytes_3453(matchBytes[3453]),
.io_matchBytes_3454(matchBytes[3454]),
.io_matchBytes_3455(matchBytes[3455]),
.io_matchBytes_3456(matchBytes[3456]),
.io_matchBytes_3457(matchBytes[3457]),
.io_matchBytes_3458(matchBytes[3458]),
.io_matchBytes_3459(matchBytes[3459]),
.io_matchBytes_3460(matchBytes[3460]),
.io_matchBytes_3461(matchBytes[3461]),
.io_matchBytes_3462(matchBytes[3462]),
.io_matchBytes_3463(matchBytes[3463]),
.io_matchBytes_3464(matchBytes[3464]),
.io_matchBytes_3465(matchBytes[3465]),
.io_matchBytes_3466(matchBytes[3466]),
.io_matchBytes_3467(matchBytes[3467]),
.io_matchBytes_3468(matchBytes[3468]),
.io_matchBytes_3469(matchBytes[3469]),
.io_matchBytes_3470(matchBytes[3470]),
.io_matchBytes_3471(matchBytes[3471]),
.io_matchBytes_3472(matchBytes[3472]),
.io_matchBytes_3473(matchBytes[3473]),
.io_matchBytes_3474(matchBytes[3474]),
.io_matchBytes_3475(matchBytes[3475]),
.io_matchBytes_3476(matchBytes[3476]),
.io_matchBytes_3477(matchBytes[3477]),
.io_matchBytes_3478(matchBytes[3478]),
.io_matchBytes_3479(matchBytes[3479]),
.io_matchBytes_3480(matchBytes[3480]),
.io_matchBytes_3481(matchBytes[3481]),
.io_matchBytes_3482(matchBytes[3482]),
.io_matchBytes_3483(matchBytes[3483]),
.io_matchBytes_3484(matchBytes[3484]),
.io_matchBytes_3485(matchBytes[3485]),
.io_matchBytes_3486(matchBytes[3486]),
.io_matchBytes_3487(matchBytes[3487]),
.io_matchBytes_3488(matchBytes[3488]),
.io_matchBytes_3489(matchBytes[3489]),
.io_matchBytes_3490(matchBytes[3490]),
.io_matchBytes_3491(matchBytes[3491]),
.io_matchBytes_3492(matchBytes[3492]),
.io_matchBytes_3493(matchBytes[3493]),
.io_matchBytes_3494(matchBytes[3494]),
.io_matchBytes_3495(matchBytes[3495]),
.io_matchBytes_3496(matchBytes[3496]),
.io_matchBytes_3497(matchBytes[3497]),
.io_matchBytes_3498(matchBytes[3498]),
.io_matchBytes_3499(matchBytes[3499]),
.io_matchBytes_3500(matchBytes[3500]),
.io_matchBytes_3501(matchBytes[3501]),
.io_matchBytes_3502(matchBytes[3502]),
.io_matchBytes_3503(matchBytes[3503]),
.io_matchBytes_3504(matchBytes[3504]),
.io_matchBytes_3505(matchBytes[3505]),
.io_matchBytes_3506(matchBytes[3506]),
.io_matchBytes_3507(matchBytes[3507]),
.io_matchBytes_3508(matchBytes[3508]),
.io_matchBytes_3509(matchBytes[3509]),
.io_matchBytes_3510(matchBytes[3510]),
.io_matchBytes_3511(matchBytes[3511]),
.io_matchBytes_3512(matchBytes[3512]),
.io_matchBytes_3513(matchBytes[3513]),
.io_matchBytes_3514(matchBytes[3514]),
.io_matchBytes_3515(matchBytes[3515]),
.io_matchBytes_3516(matchBytes[3516]),
.io_matchBytes_3517(matchBytes[3517]),
.io_matchBytes_3518(matchBytes[3518]),
.io_matchBytes_3519(matchBytes[3519]),
.io_matchBytes_3520(matchBytes[3520]),
.io_matchBytes_3521(matchBytes[3521]),
.io_matchBytes_3522(matchBytes[3522]),
.io_matchBytes_3523(matchBytes[3523]),
.io_matchBytes_3524(matchBytes[3524]),
.io_matchBytes_3525(matchBytes[3525]),
.io_matchBytes_3526(matchBytes[3526]),
.io_matchBytes_3527(matchBytes[3527]),
.io_matchBytes_3528(matchBytes[3528]),
.io_matchBytes_3529(matchBytes[3529]),
.io_matchBytes_3530(matchBytes[3530]),
.io_matchBytes_3531(matchBytes[3531]),
.io_matchBytes_3532(matchBytes[3532]),
.io_matchBytes_3533(matchBytes[3533]),
.io_matchBytes_3534(matchBytes[3534]),
.io_matchBytes_3535(matchBytes[3535]),
.io_matchBytes_3536(matchBytes[3536]),
.io_matchBytes_3537(matchBytes[3537]),
.io_matchBytes_3538(matchBytes[3538]),
.io_matchBytes_3539(matchBytes[3539]),
.io_matchBytes_3540(matchBytes[3540]),
.io_matchBytes_3541(matchBytes[3541]),
.io_matchBytes_3542(matchBytes[3542]),
.io_matchBytes_3543(matchBytes[3543]),
.io_matchBytes_3544(matchBytes[3544]),
.io_matchBytes_3545(matchBytes[3545]),
.io_matchBytes_3546(matchBytes[3546]),
.io_matchBytes_3547(matchBytes[3547]),
.io_matchBytes_3548(matchBytes[3548]),
.io_matchBytes_3549(matchBytes[3549]),
.io_matchBytes_3550(matchBytes[3550]),
.io_matchBytes_3551(matchBytes[3551]),
.io_matchBytes_3552(matchBytes[3552]),
.io_matchBytes_3553(matchBytes[3553]),
.io_matchBytes_3554(matchBytes[3554]),
.io_matchBytes_3555(matchBytes[3555]),
.io_matchBytes_3556(matchBytes[3556]),
.io_matchBytes_3557(matchBytes[3557]),
.io_matchBytes_3558(matchBytes[3558]),
.io_matchBytes_3559(matchBytes[3559]),
.io_matchBytes_3560(matchBytes[3560]),
.io_matchBytes_3561(matchBytes[3561]),
.io_matchBytes_3562(matchBytes[3562]),
.io_matchBytes_3563(matchBytes[3563]),
.io_matchBytes_3564(matchBytes[3564]),
.io_matchBytes_3565(matchBytes[3565]),
.io_matchBytes_3566(matchBytes[3566]),
.io_matchBytes_3567(matchBytes[3567]),
.io_matchBytes_3568(matchBytes[3568]),
.io_matchBytes_3569(matchBytes[3569]),
.io_matchBytes_3570(matchBytes[3570]),
.io_matchBytes_3571(matchBytes[3571]),
.io_matchBytes_3572(matchBytes[3572]),
.io_matchBytes_3573(matchBytes[3573]),
.io_matchBytes_3574(matchBytes[3574]),
.io_matchBytes_3575(matchBytes[3575]),
.io_matchBytes_3576(matchBytes[3576]),
.io_matchBytes_3577(matchBytes[3577]),
.io_matchBytes_3578(matchBytes[3578]),
.io_matchBytes_3579(matchBytes[3579]),
.io_matchBytes_3580(matchBytes[3580]),
.io_matchBytes_3581(matchBytes[3581]),
.io_matchBytes_3582(matchBytes[3582]),
.io_matchBytes_3583(matchBytes[3583]),
.io_matchBytes_3584(matchBytes[3584]),
.io_matchBytes_3585(matchBytes[3585]),
.io_matchBytes_3586(matchBytes[3586]),
.io_matchBytes_3587(matchBytes[3587]),
.io_matchBytes_3588(matchBytes[3588]),
.io_matchBytes_3589(matchBytes[3589]),
.io_matchBytes_3590(matchBytes[3590]),
.io_matchBytes_3591(matchBytes[3591]),
.io_matchBytes_3592(matchBytes[3592]),
.io_matchBytes_3593(matchBytes[3593]),
.io_matchBytes_3594(matchBytes[3594]),
.io_matchBytes_3595(matchBytes[3595]),
.io_matchBytes_3596(matchBytes[3596]),
.io_matchBytes_3597(matchBytes[3597]),
.io_matchBytes_3598(matchBytes[3598]),
.io_matchBytes_3599(matchBytes[3599]),
.io_matchBytes_3600(matchBytes[3600]),
.io_matchBytes_3601(matchBytes[3601]),
.io_matchBytes_3602(matchBytes[3602]),
.io_matchBytes_3603(matchBytes[3603]),
.io_matchBytes_3604(matchBytes[3604]),
.io_matchBytes_3605(matchBytes[3605]),
.io_matchBytes_3606(matchBytes[3606]),
.io_matchBytes_3607(matchBytes[3607]),
.io_matchBytes_3608(matchBytes[3608]),
.io_matchBytes_3609(matchBytes[3609]),
.io_matchBytes_3610(matchBytes[3610]),
.io_matchBytes_3611(matchBytes[3611]),
.io_matchBytes_3612(matchBytes[3612]),
.io_matchBytes_3613(matchBytes[3613]),
.io_matchBytes_3614(matchBytes[3614]),
.io_matchBytes_3615(matchBytes[3615]),
.io_matchBytes_3616(matchBytes[3616]),
.io_matchBytes_3617(matchBytes[3617]),
.io_matchBytes_3618(matchBytes[3618]),
.io_matchBytes_3619(matchBytes[3619]),
.io_matchBytes_3620(matchBytes[3620]),
.io_matchBytes_3621(matchBytes[3621]),
.io_matchBytes_3622(matchBytes[3622]),
.io_matchBytes_3623(matchBytes[3623]),
.io_matchBytes_3624(matchBytes[3624]),
.io_matchBytes_3625(matchBytes[3625]),
.io_matchBytes_3626(matchBytes[3626]),
.io_matchBytes_3627(matchBytes[3627]),
.io_matchBytes_3628(matchBytes[3628]),
.io_matchBytes_3629(matchBytes[3629]),
.io_matchBytes_3630(matchBytes[3630]),
.io_matchBytes_3631(matchBytes[3631]),
.io_matchBytes_3632(matchBytes[3632]),
.io_matchBytes_3633(matchBytes[3633]),
.io_matchBytes_3634(matchBytes[3634]),
.io_matchBytes_3635(matchBytes[3635]),
.io_matchBytes_3636(matchBytes[3636]),
.io_matchBytes_3637(matchBytes[3637]),
.io_matchBytes_3638(matchBytes[3638]),
.io_matchBytes_3639(matchBytes[3639]),
.io_matchBytes_3640(matchBytes[3640]),
.io_matchBytes_3641(matchBytes[3641]),
.io_matchBytes_3642(matchBytes[3642]),
.io_matchBytes_3643(matchBytes[3643]),
.io_matchBytes_3644(matchBytes[3644]),
.io_matchBytes_3645(matchBytes[3645]),
.io_matchBytes_3646(matchBytes[3646]),
.io_matchBytes_3647(matchBytes[3647]),
.io_matchBytes_3648(matchBytes[3648]),
.io_matchBytes_3649(matchBytes[3649]),
.io_matchBytes_3650(matchBytes[3650]),
.io_matchBytes_3651(matchBytes[3651]),
.io_matchBytes_3652(matchBytes[3652]),
.io_matchBytes_3653(matchBytes[3653]),
.io_matchBytes_3654(matchBytes[3654]),
.io_matchBytes_3655(matchBytes[3655]),
.io_matchBytes_3656(matchBytes[3656]),
.io_matchBytes_3657(matchBytes[3657]),
.io_matchBytes_3658(matchBytes[3658]),
.io_matchBytes_3659(matchBytes[3659]),
.io_matchBytes_3660(matchBytes[3660]),
.io_matchBytes_3661(matchBytes[3661]),
.io_matchBytes_3662(matchBytes[3662]),
.io_matchBytes_3663(matchBytes[3663]),
.io_matchBytes_3664(matchBytes[3664]),
.io_matchBytes_3665(matchBytes[3665]),
.io_matchBytes_3666(matchBytes[3666]),
.io_matchBytes_3667(matchBytes[3667]),
.io_matchBytes_3668(matchBytes[3668]),
.io_matchBytes_3669(matchBytes[3669]),
.io_matchBytes_3670(matchBytes[3670]),
.io_matchBytes_3671(matchBytes[3671]),
.io_matchBytes_3672(matchBytes[3672]),
.io_matchBytes_3673(matchBytes[3673]),
.io_matchBytes_3674(matchBytes[3674]),
.io_matchBytes_3675(matchBytes[3675]),
.io_matchBytes_3676(matchBytes[3676]),
.io_matchBytes_3677(matchBytes[3677]),
.io_matchBytes_3678(matchBytes[3678]),
.io_matchBytes_3679(matchBytes[3679]),
.io_matchBytes_3680(matchBytes[3680]),
.io_matchBytes_3681(matchBytes[3681]),
.io_matchBytes_3682(matchBytes[3682]),
.io_matchBytes_3683(matchBytes[3683]),
.io_matchBytes_3684(matchBytes[3684]),
.io_matchBytes_3685(matchBytes[3685]),
.io_matchBytes_3686(matchBytes[3686]),
.io_matchBytes_3687(matchBytes[3687]),
.io_matchBytes_3688(matchBytes[3688]),
.io_matchBytes_3689(matchBytes[3689]),
.io_matchBytes_3690(matchBytes[3690]),
.io_matchBytes_3691(matchBytes[3691]),
.io_matchBytes_3692(matchBytes[3692]),
.io_matchBytes_3693(matchBytes[3693]),
.io_matchBytes_3694(matchBytes[3694]),
.io_matchBytes_3695(matchBytes[3695]),
.io_matchBytes_3696(matchBytes[3696]),
.io_matchBytes_3697(matchBytes[3697]),
.io_matchBytes_3698(matchBytes[3698]),
.io_matchBytes_3699(matchBytes[3699]),
.io_matchBytes_3700(matchBytes[3700]),
.io_matchBytes_3701(matchBytes[3701]),
.io_matchBytes_3702(matchBytes[3702]),
.io_matchBytes_3703(matchBytes[3703]),
.io_matchBytes_3704(matchBytes[3704]),
.io_matchBytes_3705(matchBytes[3705]),
.io_matchBytes_3706(matchBytes[3706]),
.io_matchBytes_3707(matchBytes[3707]),
.io_matchBytes_3708(matchBytes[3708]),
.io_matchBytes_3709(matchBytes[3709]),
.io_matchBytes_3710(matchBytes[3710]),
.io_matchBytes_3711(matchBytes[3711]),
.io_matchBytes_3712(matchBytes[3712]),
.io_matchBytes_3713(matchBytes[3713]),
.io_matchBytes_3714(matchBytes[3714]),
.io_matchBytes_3715(matchBytes[3715]),
.io_matchBytes_3716(matchBytes[3716]),
.io_matchBytes_3717(matchBytes[3717]),
.io_matchBytes_3718(matchBytes[3718]),
.io_matchBytes_3719(matchBytes[3719]),
.io_matchBytes_3720(matchBytes[3720]),
.io_matchBytes_3721(matchBytes[3721]),
.io_matchBytes_3722(matchBytes[3722]),
.io_matchBytes_3723(matchBytes[3723]),
.io_matchBytes_3724(matchBytes[3724]),
.io_matchBytes_3725(matchBytes[3725]),
.io_matchBytes_3726(matchBytes[3726]),
.io_matchBytes_3727(matchBytes[3727]),
.io_matchBytes_3728(matchBytes[3728]),
.io_matchBytes_3729(matchBytes[3729]),
.io_matchBytes_3730(matchBytes[3730]),
.io_matchBytes_3731(matchBytes[3731]),
.io_matchBytes_3732(matchBytes[3732]),
.io_matchBytes_3733(matchBytes[3733]),
.io_matchBytes_3734(matchBytes[3734]),
.io_matchBytes_3735(matchBytes[3735]),
.io_matchBytes_3736(matchBytes[3736]),
.io_matchBytes_3737(matchBytes[3737]),
.io_matchBytes_3738(matchBytes[3738]),
.io_matchBytes_3739(matchBytes[3739]),
.io_matchBytes_3740(matchBytes[3740]),
.io_matchBytes_3741(matchBytes[3741]),
.io_matchBytes_3742(matchBytes[3742]),
.io_matchBytes_3743(matchBytes[3743]),
.io_matchBytes_3744(matchBytes[3744]),
.io_matchBytes_3745(matchBytes[3745]),
.io_matchBytes_3746(matchBytes[3746]),
.io_matchBytes_3747(matchBytes[3747]),
.io_matchBytes_3748(matchBytes[3748]),
.io_matchBytes_3749(matchBytes[3749]),
.io_matchBytes_3750(matchBytes[3750]),
.io_matchBytes_3751(matchBytes[3751]),
.io_matchBytes_3752(matchBytes[3752]),
.io_matchBytes_3753(matchBytes[3753]),
.io_matchBytes_3754(matchBytes[3754]),
.io_matchBytes_3755(matchBytes[3755]),
.io_matchBytes_3756(matchBytes[3756]),
.io_matchBytes_3757(matchBytes[3757]),
.io_matchBytes_3758(matchBytes[3758]),
.io_matchBytes_3759(matchBytes[3759]),
.io_matchBytes_3760(matchBytes[3760]),
.io_matchBytes_3761(matchBytes[3761]),
.io_matchBytes_3762(matchBytes[3762]),
.io_matchBytes_3763(matchBytes[3763]),
.io_matchBytes_3764(matchBytes[3764]),
.io_matchBytes_3765(matchBytes[3765]),
.io_matchBytes_3766(matchBytes[3766]),
.io_matchBytes_3767(matchBytes[3767]),
.io_matchBytes_3768(matchBytes[3768]),
.io_matchBytes_3769(matchBytes[3769]),
.io_matchBytes_3770(matchBytes[3770]),
.io_matchBytes_3771(matchBytes[3771]),
.io_matchBytes_3772(matchBytes[3772]),
.io_matchBytes_3773(matchBytes[3773]),
.io_matchBytes_3774(matchBytes[3774]),
.io_matchBytes_3775(matchBytes[3775]),
.io_matchBytes_3776(matchBytes[3776]),
.io_matchBytes_3777(matchBytes[3777]),
.io_matchBytes_3778(matchBytes[3778]),
.io_matchBytes_3779(matchBytes[3779]),
.io_matchBytes_3780(matchBytes[3780]),
.io_matchBytes_3781(matchBytes[3781]),
.io_matchBytes_3782(matchBytes[3782]),
.io_matchBytes_3783(matchBytes[3783]),
.io_matchBytes_3784(matchBytes[3784]),
.io_matchBytes_3785(matchBytes[3785]),
.io_matchBytes_3786(matchBytes[3786]),
.io_matchBytes_3787(matchBytes[3787]),
.io_matchBytes_3788(matchBytes[3788]),
.io_matchBytes_3789(matchBytes[3789]),
.io_matchBytes_3790(matchBytes[3790]),
.io_matchBytes_3791(matchBytes[3791]),
.io_matchBytes_3792(matchBytes[3792]),
.io_matchBytes_3793(matchBytes[3793]),
.io_matchBytes_3794(matchBytes[3794]),
.io_matchBytes_3795(matchBytes[3795]),
.io_matchBytes_3796(matchBytes[3796]),
.io_matchBytes_3797(matchBytes[3797]),
.io_matchBytes_3798(matchBytes[3798]),
.io_matchBytes_3799(matchBytes[3799]),
.io_matchBytes_3800(matchBytes[3800]),
.io_matchBytes_3801(matchBytes[3801]),
.io_matchBytes_3802(matchBytes[3802]),
.io_matchBytes_3803(matchBytes[3803]),
.io_matchBytes_3804(matchBytes[3804]),
.io_matchBytes_3805(matchBytes[3805]),
.io_matchBytes_3806(matchBytes[3806]),
.io_matchBytes_3807(matchBytes[3807]),
.io_matchBytes_3808(matchBytes[3808]),
.io_matchBytes_3809(matchBytes[3809]),
.io_matchBytes_3810(matchBytes[3810]),
.io_matchBytes_3811(matchBytes[3811]),
.io_matchBytes_3812(matchBytes[3812]),
.io_matchBytes_3813(matchBytes[3813]),
.io_matchBytes_3814(matchBytes[3814]),
.io_matchBytes_3815(matchBytes[3815]),
.io_matchBytes_3816(matchBytes[3816]),
.io_matchBytes_3817(matchBytes[3817]),
.io_matchBytes_3818(matchBytes[3818]),
.io_matchBytes_3819(matchBytes[3819]),
.io_matchBytes_3820(matchBytes[3820]),
.io_matchBytes_3821(matchBytes[3821]),
.io_matchBytes_3822(matchBytes[3822]),
.io_matchBytes_3823(matchBytes[3823]),
.io_matchBytes_3824(matchBytes[3824]),
.io_matchBytes_3825(matchBytes[3825]),
.io_matchBytes_3826(matchBytes[3826]),
.io_matchBytes_3827(matchBytes[3827]),
.io_matchBytes_3828(matchBytes[3828]),
.io_matchBytes_3829(matchBytes[3829]),
.io_matchBytes_3830(matchBytes[3830]),
.io_matchBytes_3831(matchBytes[3831]),
.io_matchBytes_3832(matchBytes[3832]),
.io_matchBytes_3833(matchBytes[3833]),
.io_matchBytes_3834(matchBytes[3834]),
.io_matchBytes_3835(matchBytes[3835]),
.io_matchBytes_3836(matchBytes[3836]),
.io_matchBytes_3837(matchBytes[3837]),
.io_matchBytes_3838(matchBytes[3838]),
.io_matchBytes_3839(matchBytes[3839]),
.io_matchBytes_3840(matchBytes[3840]),
.io_matchBytes_3841(matchBytes[3841]),
.io_matchBytes_3842(matchBytes[3842]),
.io_matchBytes_3843(matchBytes[3843]),
.io_matchBytes_3844(matchBytes[3844]),
.io_matchBytes_3845(matchBytes[3845]),
.io_matchBytes_3846(matchBytes[3846]),
.io_matchBytes_3847(matchBytes[3847]),
.io_matchBytes_3848(matchBytes[3848]),
.io_matchBytes_3849(matchBytes[3849]),
.io_matchBytes_3850(matchBytes[3850]),
.io_matchBytes_3851(matchBytes[3851]),
.io_matchBytes_3852(matchBytes[3852]),
.io_matchBytes_3853(matchBytes[3853]),
.io_matchBytes_3854(matchBytes[3854]),
.io_matchBytes_3855(matchBytes[3855]),
.io_matchBytes_3856(matchBytes[3856]),
.io_matchBytes_3857(matchBytes[3857]),
.io_matchBytes_3858(matchBytes[3858]),
.io_matchBytes_3859(matchBytes[3859]),
.io_matchBytes_3860(matchBytes[3860]),
.io_matchBytes_3861(matchBytes[3861]),
.io_matchBytes_3862(matchBytes[3862]),
.io_matchBytes_3863(matchBytes[3863]),
.io_matchBytes_3864(matchBytes[3864]),
.io_matchBytes_3865(matchBytes[3865]),
.io_matchBytes_3866(matchBytes[3866]),
.io_matchBytes_3867(matchBytes[3867]),
.io_matchBytes_3868(matchBytes[3868]),
.io_matchBytes_3869(matchBytes[3869]),
.io_matchBytes_3870(matchBytes[3870]),
.io_matchBytes_3871(matchBytes[3871]),
.io_matchBytes_3872(matchBytes[3872]),
.io_matchBytes_3873(matchBytes[3873]),
.io_matchBytes_3874(matchBytes[3874]),
.io_matchBytes_3875(matchBytes[3875]),
.io_matchBytes_3876(matchBytes[3876]),
.io_matchBytes_3877(matchBytes[3877]),
.io_matchBytes_3878(matchBytes[3878]),
.io_matchBytes_3879(matchBytes[3879]),
.io_matchBytes_3880(matchBytes[3880]),
.io_matchBytes_3881(matchBytes[3881]),
.io_matchBytes_3882(matchBytes[3882]),
.io_matchBytes_3883(matchBytes[3883]),
.io_matchBytes_3884(matchBytes[3884]),
.io_matchBytes_3885(matchBytes[3885]),
.io_matchBytes_3886(matchBytes[3886]),
.io_matchBytes_3887(matchBytes[3887]),
.io_matchBytes_3888(matchBytes[3888]),
.io_matchBytes_3889(matchBytes[3889]),
.io_matchBytes_3890(matchBytes[3890]),
.io_matchBytes_3891(matchBytes[3891]),
.io_matchBytes_3892(matchBytes[3892]),
.io_matchBytes_3893(matchBytes[3893]),
.io_matchBytes_3894(matchBytes[3894]),
.io_matchBytes_3895(matchBytes[3895]),
.io_matchBytes_3896(matchBytes[3896]),
.io_matchBytes_3897(matchBytes[3897]),
.io_matchBytes_3898(matchBytes[3898]),
.io_matchBytes_3899(matchBytes[3899]),
.io_matchBytes_3900(matchBytes[3900]),
.io_matchBytes_3901(matchBytes[3901]),
.io_matchBytes_3902(matchBytes[3902]),
.io_matchBytes_3903(matchBytes[3903]),
.io_matchBytes_3904(matchBytes[3904]),
.io_matchBytes_3905(matchBytes[3905]),
.io_matchBytes_3906(matchBytes[3906]),
.io_matchBytes_3907(matchBytes[3907]),
.io_matchBytes_3908(matchBytes[3908]),
.io_matchBytes_3909(matchBytes[3909]),
.io_matchBytes_3910(matchBytes[3910]),
.io_matchBytes_3911(matchBytes[3911]),
.io_matchBytes_3912(matchBytes[3912]),
.io_matchBytes_3913(matchBytes[3913]),
.io_matchBytes_3914(matchBytes[3914]),
.io_matchBytes_3915(matchBytes[3915]),
.io_matchBytes_3916(matchBytes[3916]),
.io_matchBytes_3917(matchBytes[3917]),
.io_matchBytes_3918(matchBytes[3918]),
.io_matchBytes_3919(matchBytes[3919]),
.io_matchBytes_3920(matchBytes[3920]),
.io_matchBytes_3921(matchBytes[3921]),
.io_matchBytes_3922(matchBytes[3922]),
.io_matchBytes_3923(matchBytes[3923]),
.io_matchBytes_3924(matchBytes[3924]),
.io_matchBytes_3925(matchBytes[3925]),
.io_matchBytes_3926(matchBytes[3926]),
.io_matchBytes_3927(matchBytes[3927]),
.io_matchBytes_3928(matchBytes[3928]),
.io_matchBytes_3929(matchBytes[3929]),
.io_matchBytes_3930(matchBytes[3930]),
.io_matchBytes_3931(matchBytes[3931]),
.io_matchBytes_3932(matchBytes[3932]),
.io_matchBytes_3933(matchBytes[3933]),
.io_matchBytes_3934(matchBytes[3934]),
.io_matchBytes_3935(matchBytes[3935]),
.io_matchBytes_3936(matchBytes[3936]),
.io_matchBytes_3937(matchBytes[3937]),
.io_matchBytes_3938(matchBytes[3938]),
.io_matchBytes_3939(matchBytes[3939]),
.io_matchBytes_3940(matchBytes[3940]),
.io_matchBytes_3941(matchBytes[3941]),
.io_matchBytes_3942(matchBytes[3942]),
.io_matchBytes_3943(matchBytes[3943]),
.io_matchBytes_3944(matchBytes[3944]),
.io_matchBytes_3945(matchBytes[3945]),
.io_matchBytes_3946(matchBytes[3946]),
.io_matchBytes_3947(matchBytes[3947]),
.io_matchBytes_3948(matchBytes[3948]),
.io_matchBytes_3949(matchBytes[3949]),
.io_matchBytes_3950(matchBytes[3950]),
.io_matchBytes_3951(matchBytes[3951]),
.io_matchBytes_3952(matchBytes[3952]),
.io_matchBytes_3953(matchBytes[3953]),
.io_matchBytes_3954(matchBytes[3954]),
.io_matchBytes_3955(matchBytes[3955]),
.io_matchBytes_3956(matchBytes[3956]),
.io_matchBytes_3957(matchBytes[3957]),
.io_matchBytes_3958(matchBytes[3958]),
.io_matchBytes_3959(matchBytes[3959]),
.io_matchBytes_3960(matchBytes[3960]),
.io_matchBytes_3961(matchBytes[3961]),
.io_matchBytes_3962(matchBytes[3962]),
.io_matchBytes_3963(matchBytes[3963]),
.io_matchBytes_3964(matchBytes[3964]),
.io_matchBytes_3965(matchBytes[3965]),
.io_matchBytes_3966(matchBytes[3966]),
.io_matchBytes_3967(matchBytes[3967]),
.io_matchBytes_3968(matchBytes[3968]),
.io_matchBytes_3969(matchBytes[3969]),
.io_matchBytes_3970(matchBytes[3970]),
.io_matchBytes_3971(matchBytes[3971]),
.io_matchBytes_3972(matchBytes[3972]),
.io_matchBytes_3973(matchBytes[3973]),
.io_matchBytes_3974(matchBytes[3974]),
.io_matchBytes_3975(matchBytes[3975]),
.io_matchBytes_3976(matchBytes[3976]),
.io_matchBytes_3977(matchBytes[3977]),
.io_matchBytes_3978(matchBytes[3978]),
.io_matchBytes_3979(matchBytes[3979]),
.io_matchBytes_3980(matchBytes[3980]),
.io_matchBytes_3981(matchBytes[3981]),
.io_matchBytes_3982(matchBytes[3982]),
.io_matchBytes_3983(matchBytes[3983]),
.io_matchBytes_3984(matchBytes[3984]),
.io_matchBytes_3985(matchBytes[3985]),
.io_matchBytes_3986(matchBytes[3986]),
.io_matchBytes_3987(matchBytes[3987]),
.io_matchBytes_3988(matchBytes[3988]),
.io_matchBytes_3989(matchBytes[3989]),
.io_matchBytes_3990(matchBytes[3990]),
.io_matchBytes_3991(matchBytes[3991]),
.io_matchBytes_3992(matchBytes[3992]),
.io_matchBytes_3993(matchBytes[3993]),
.io_matchBytes_3994(matchBytes[3994]),
.io_matchBytes_3995(matchBytes[3995]),
.io_matchBytes_3996(matchBytes[3996]),
.io_matchBytes_3997(matchBytes[3997]),
.io_matchBytes_3998(matchBytes[3998]),
.io_matchBytes_3999(matchBytes[3999]),
.io_matchBytes_4000(matchBytes[4000]),
.io_matchBytes_4001(matchBytes[4001]),
.io_matchBytes_4002(matchBytes[4002]),
.io_matchBytes_4003(matchBytes[4003]),
.io_matchBytes_4004(matchBytes[4004]),
.io_matchBytes_4005(matchBytes[4005]),
.io_matchBytes_4006(matchBytes[4006]),
.io_matchBytes_4007(matchBytes[4007]),
.io_matchBytes_4008(matchBytes[4008]),
.io_matchBytes_4009(matchBytes[4009]),
.io_matchBytes_4010(matchBytes[4010]),
.io_matchBytes_4011(matchBytes[4011]),
.io_matchBytes_4012(matchBytes[4012]),
.io_matchBytes_4013(matchBytes[4013]),
.io_matchBytes_4014(matchBytes[4014]),
.io_matchBytes_4015(matchBytes[4015]),
.io_matchBytes_4016(matchBytes[4016]),
.io_matchBytes_4017(matchBytes[4017]),
.io_matchBytes_4018(matchBytes[4018]),
.io_matchBytes_4019(matchBytes[4019]),
.io_matchBytes_4020(matchBytes[4020]),
.io_matchBytes_4021(matchBytes[4021]),
.io_matchBytes_4022(matchBytes[4022]),
.io_matchBytes_4023(matchBytes[4023]),
.io_matchBytes_4024(matchBytes[4024]),
.io_matchBytes_4025(matchBytes[4025]),
.io_matchBytes_4026(matchBytes[4026]),
.io_matchBytes_4027(matchBytes[4027]),
.io_matchBytes_4028(matchBytes[4028]),
.io_matchBytes_4029(matchBytes[4029]),
.io_matchBytes_4030(matchBytes[4030]),
.io_matchBytes_4031(matchBytes[4031]),
.io_matchBytes_4032(matchBytes[4032]),
.io_matchBytes_4033(matchBytes[4033]),
.io_matchBytes_4034(matchBytes[4034]),
.io_matchBytes_4035(matchBytes[4035]),
.io_matchBytes_4036(matchBytes[4036]),
.io_matchBytes_4037(matchBytes[4037]),
.io_matchBytes_4038(matchBytes[4038]),
.io_matchBytes_4039(matchBytes[4039]),
.io_matchBytes_4040(matchBytes[4040]),
.io_matchBytes_4041(matchBytes[4041]),
.io_matchBytes_4042(matchBytes[4042]),
.io_matchBytes_4043(matchBytes[4043]),
.io_matchBytes_4044(matchBytes[4044]),
.io_matchBytes_4045(matchBytes[4045]),
.io_matchBytes_4046(matchBytes[4046]),
.io_matchBytes_4047(matchBytes[4047]),
.io_matchBytes_4048(matchBytes[4048]),
.io_matchBytes_4049(matchBytes[4049]),
.io_matchBytes_4050(matchBytes[4050]),
.io_matchBytes_4051(matchBytes[4051]),
.io_matchBytes_4052(matchBytes[4052]),
.io_matchBytes_4053(matchBytes[4053]),
.io_matchBytes_4054(matchBytes[4054]),
.io_matchBytes_4055(matchBytes[4055]),
.io_matchBytes_4056(matchBytes[4056]),
.io_matchBytes_4057(matchBytes[4057]),
.io_matchBytes_4058(matchBytes[4058]),
.io_matchBytes_4059(matchBytes[4059]),
.io_matchBytes_4060(matchBytes[4060]),
.io_matchBytes_4061(matchBytes[4061]),
.io_matchBytes_4062(matchBytes[4062]),
.io_matchBytes_4063(matchBytes[4063]),
.io_matchBytes_4064(matchBytes[4064]),
.io_matchBytes_4065(matchBytes[4065]),
.io_matchBytes_4066(matchBytes[4066]),
.io_matchBytes_4067(matchBytes[4067]),
.io_matchBytes_4068(matchBytes[4068]),
.io_matchBytes_4069(matchBytes[4069]),
.io_matchBytes_4070(matchBytes[4070]),
.io_matchBytes_4071(matchBytes[4071]),
.io_matchBytes_4072(matchBytes[4072]),
.io_matchBytes_4073(matchBytes[4073]),
.io_matchBytes_4074(matchBytes[4074]),
.io_matchBytes_4075(matchBytes[4075]),
.io_matchBytes_4076(matchBytes[4076]),
.io_matchBytes_4077(matchBytes[4077]),
.io_matchBytes_4078(matchBytes[4078]),
.io_matchBytes_4079(matchBytes[4079]),
.io_matchBytes_4080(matchBytes[4080]),
.io_matchBytes_4081(matchBytes[4081]),
.io_matchBytes_4082(matchBytes[4082]),
.io_matchBytes_4083(matchBytes[4083]),
.io_matchBytes_4084(matchBytes[4084]),
.io_matchBytes_4085(matchBytes[4085]),
.io_matchBytes_4086(matchBytes[4086]),
.io_matchBytes_4087(matchBytes[4087]),
.io_matchBytes_4088(matchBytes[4088]),
.io_matchBytes_4089(matchBytes[4089]),
.io_matchBytes_4090(matchBytes[4090]),
.io_matchBytes_4091(matchBytes[4091]),
.io_matchBytes_4092(matchBytes[4092]),
.io_matchBytes_4093(matchBytes[4093]),
.io_matchBytes_4094(matchBytes[4094]),
.io_matchBytes_4095(matchBytes[4095]),
.io_completeMatch(completeMatch),
.io_outputBytes(outputBytes),
.io_finished(finished)
         );

endmodule

